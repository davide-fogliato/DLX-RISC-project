
module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n33, n66, n67, n100;

  BUF_X1 U1 ( .A(n100), .Z(n33) );
  BUF_X1 U2 ( .A(n100), .Z(n66) );
  BUF_X1 U3 ( .A(n100), .Z(n67) );
  INV_X1 U4 ( .A(n62), .ZN(Y[12]) );
  AOI22_X1 U5 ( .A1(A[12]), .A2(n33), .B1(B[12]), .B2(SEL), .ZN(n62) );
  INV_X1 U6 ( .A(n61), .ZN(Y[13]) );
  AOI22_X1 U7 ( .A1(A[13]), .A2(n33), .B1(B[13]), .B2(SEL), .ZN(n61) );
  INV_X1 U8 ( .A(n59), .ZN(Y[15]) );
  AOI22_X1 U9 ( .A1(A[15]), .A2(n33), .B1(B[15]), .B2(SEL), .ZN(n59) );
  INV_X1 U10 ( .A(n58), .ZN(Y[16]) );
  AOI22_X1 U11 ( .A1(A[16]), .A2(n33), .B1(B[16]), .B2(SEL), .ZN(n58) );
  INV_X1 U12 ( .A(n56), .ZN(Y[18]) );
  AOI22_X1 U13 ( .A1(A[18]), .A2(n33), .B1(B[18]), .B2(SEL), .ZN(n56) );
  INV_X1 U14 ( .A(n55), .ZN(Y[19]) );
  AOI22_X1 U15 ( .A1(A[19]), .A2(n33), .B1(B[19]), .B2(SEL), .ZN(n55) );
  INV_X1 U16 ( .A(n53), .ZN(Y[20]) );
  AOI22_X1 U17 ( .A1(A[20]), .A2(n66), .B1(B[20]), .B2(SEL), .ZN(n53) );
  INV_X1 U18 ( .A(n51), .ZN(Y[22]) );
  AOI22_X1 U19 ( .A1(A[22]), .A2(n66), .B1(B[22]), .B2(SEL), .ZN(n51) );
  INV_X1 U20 ( .A(n50), .ZN(Y[23]) );
  AOI22_X1 U21 ( .A1(A[23]), .A2(n66), .B1(B[23]), .B2(SEL), .ZN(n50) );
  INV_X1 U22 ( .A(n49), .ZN(Y[24]) );
  AOI22_X1 U23 ( .A1(A[24]), .A2(n66), .B1(B[24]), .B2(SEL), .ZN(n49) );
  INV_X1 U24 ( .A(n48), .ZN(Y[25]) );
  AOI22_X1 U25 ( .A1(A[25]), .A2(n66), .B1(B[25]), .B2(SEL), .ZN(n48) );
  INV_X1 U26 ( .A(n47), .ZN(Y[26]) );
  AOI22_X1 U27 ( .A1(A[26]), .A2(n66), .B1(B[26]), .B2(SEL), .ZN(n47) );
  INV_X1 U28 ( .A(n46), .ZN(Y[27]) );
  AOI22_X1 U29 ( .A1(A[27]), .A2(n66), .B1(B[27]), .B2(SEL), .ZN(n46) );
  INV_X1 U30 ( .A(n45), .ZN(Y[28]) );
  AOI22_X1 U31 ( .A1(A[28]), .A2(n66), .B1(B[28]), .B2(SEL), .ZN(n45) );
  INV_X1 U32 ( .A(n44), .ZN(Y[29]) );
  AOI22_X1 U33 ( .A1(A[29]), .A2(n66), .B1(B[29]), .B2(SEL), .ZN(n44) );
  INV_X1 U34 ( .A(n42), .ZN(Y[30]) );
  AOI22_X1 U35 ( .A1(A[30]), .A2(n66), .B1(B[30]), .B2(SEL), .ZN(n42) );
  INV_X1 U36 ( .A(n41), .ZN(Y[31]) );
  AOI22_X1 U37 ( .A1(A[31]), .A2(n67), .B1(B[31]), .B2(SEL), .ZN(n41) );
  INV_X1 U38 ( .A(n60), .ZN(Y[14]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n33), .B1(B[14]), .B2(SEL), .ZN(n60) );
  INV_X1 U40 ( .A(n57), .ZN(Y[17]) );
  AOI22_X1 U41 ( .A1(A[17]), .A2(n33), .B1(B[17]), .B2(SEL), .ZN(n57) );
  INV_X1 U42 ( .A(n52), .ZN(Y[21]) );
  AOI22_X1 U43 ( .A1(A[21]), .A2(n66), .B1(B[21]), .B2(SEL), .ZN(n52) );
  INV_X1 U44 ( .A(n36), .ZN(Y[7]) );
  AOI22_X1 U45 ( .A1(A[7]), .A2(n67), .B1(B[7]), .B2(SEL), .ZN(n36) );
  INV_X1 U46 ( .A(n40), .ZN(Y[3]) );
  AOI22_X1 U47 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(SEL), .ZN(n40) );
  INV_X1 U48 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U49 ( .A1(A[0]), .A2(n33), .B1(B[0]), .B2(SEL), .ZN(n65) );
  INV_X1 U50 ( .A(n54), .ZN(Y[1]) );
  AOI22_X1 U51 ( .A1(A[1]), .A2(n33), .B1(B[1]), .B2(SEL), .ZN(n54) );
  INV_X1 U52 ( .A(n43), .ZN(Y[2]) );
  AOI22_X1 U53 ( .A1(A[2]), .A2(n66), .B1(B[2]), .B2(SEL), .ZN(n43) );
  INV_X1 U54 ( .A(n39), .ZN(Y[4]) );
  AOI22_X1 U55 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(SEL), .ZN(n39) );
  INV_X1 U56 ( .A(n38), .ZN(Y[5]) );
  AOI22_X1 U57 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(SEL), .ZN(n38) );
  INV_X1 U58 ( .A(n37), .ZN(Y[6]) );
  AOI22_X1 U59 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(SEL), .ZN(n37) );
  INV_X1 U60 ( .A(n35), .ZN(Y[8]) );
  AOI22_X1 U61 ( .A1(A[8]), .A2(n67), .B1(B[8]), .B2(SEL), .ZN(n35) );
  INV_X1 U62 ( .A(n64), .ZN(Y[10]) );
  AOI22_X1 U63 ( .A1(A[10]), .A2(n33), .B1(B[10]), .B2(SEL), .ZN(n64) );
  INV_X1 U64 ( .A(n63), .ZN(Y[11]) );
  AOI22_X1 U65 ( .A1(A[11]), .A2(n33), .B1(B[11]), .B2(SEL), .ZN(n63) );
  INV_X1 U66 ( .A(n34), .ZN(Y[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n67), .B1(SEL), .B2(B[9]), .ZN(n34) );
  INV_X1 U68 ( .A(SEL), .ZN(n100) );
endmodule


module REG_GEN_NBIT32_0 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n47), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n47), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n47), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n47), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n47), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n47), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n47), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n47), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n47), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n47), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n47), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n47), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n48), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n48), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n48), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n48), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n48), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n48), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n48), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n48), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n48), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n48), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n48), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n48), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n49), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n49), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n49), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n49), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n49), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n49), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n49), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n49), .Q(Q[0]), .QN(n97) );
  BUF_X1 U2 ( .A(RESET_n), .Z(n48) );
  BUF_X1 U3 ( .A(RESET_n), .Z(n47) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n49) );
  INV_X1 U5 ( .A(n46), .ZN(n37) );
  INV_X1 U6 ( .A(n46), .ZN(n36) );
  BUF_X1 U7 ( .A(n35), .Z(n46) );
  BUF_X1 U8 ( .A(n34), .Z(n41) );
  BUF_X1 U9 ( .A(n34), .Z(n42) );
  BUF_X1 U10 ( .A(n35), .Z(n44) );
  BUF_X1 U11 ( .A(n33), .Z(n38) );
  BUF_X1 U12 ( .A(n33), .Z(n39) );
  BUF_X1 U13 ( .A(n33), .Z(n40) );
  BUF_X1 U14 ( .A(n34), .Z(n43) );
  BUF_X1 U15 ( .A(n35), .Z(n45) );
  OAI22_X1 U16 ( .A1(n85), .A2(n37), .B1(n42), .B2(n57), .ZN(n20) );
  INV_X1 U17 ( .A(D[12]), .ZN(n57) );
  OAI22_X1 U18 ( .A1(n84), .A2(n36), .B1(n43), .B2(n56), .ZN(n19) );
  INV_X1 U19 ( .A(D[13]), .ZN(n56) );
  OAI22_X1 U20 ( .A1(n82), .A2(n36), .B1(n43), .B2(n54), .ZN(n17) );
  INV_X1 U21 ( .A(D[15]), .ZN(n54) );
  OAI22_X1 U22 ( .A1(n81), .A2(n36), .B1(n44), .B2(n61), .ZN(n16) );
  INV_X1 U23 ( .A(D[16]), .ZN(n61) );
  OAI22_X1 U24 ( .A1(n79), .A2(n36), .B1(n44), .B2(n59), .ZN(n14) );
  INV_X1 U25 ( .A(D[18]), .ZN(n59) );
  OAI22_X1 U26 ( .A1(n78), .A2(n36), .B1(n44), .B2(n58), .ZN(n13) );
  INV_X1 U27 ( .A(D[19]), .ZN(n58) );
  OAI22_X1 U28 ( .A1(n77), .A2(n36), .B1(n45), .B2(n65), .ZN(n12) );
  INV_X1 U29 ( .A(D[20]), .ZN(n65) );
  OAI22_X1 U30 ( .A1(n75), .A2(n36), .B1(n45), .B2(n63), .ZN(n10) );
  INV_X1 U31 ( .A(D[22]), .ZN(n63) );
  OAI22_X1 U32 ( .A1(n74), .A2(n37), .B1(n38), .B2(n62), .ZN(n9) );
  INV_X1 U33 ( .A(D[23]), .ZN(n62) );
  OAI22_X1 U34 ( .A1(n73), .A2(n36), .B1(n38), .B2(n101), .ZN(n8) );
  INV_X1 U35 ( .A(D[24]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n72), .A2(n37), .B1(n38), .B2(n100), .ZN(n7) );
  INV_X1 U37 ( .A(D[25]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n71), .A2(n36), .B1(n38), .B2(n99), .ZN(n6) );
  INV_X1 U39 ( .A(D[26]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n70), .A2(n37), .B1(n39), .B2(n98), .ZN(n5) );
  INV_X1 U41 ( .A(D[27]), .ZN(n98) );
  OAI22_X1 U42 ( .A1(n69), .A2(n36), .B1(n39), .B2(n105), .ZN(n4) );
  INV_X1 U43 ( .A(D[28]), .ZN(n105) );
  OAI22_X1 U44 ( .A1(n68), .A2(n37), .B1(n40), .B2(n104), .ZN(n3) );
  INV_X1 U45 ( .A(D[29]), .ZN(n104) );
  OAI22_X1 U46 ( .A1(n67), .A2(n36), .B1(n43), .B2(n103), .ZN(n2) );
  INV_X1 U47 ( .A(D[30]), .ZN(n103) );
  OAI22_X1 U48 ( .A1(n66), .A2(n36), .B1(n45), .B2(n102), .ZN(n1) );
  INV_X1 U49 ( .A(D[31]), .ZN(n102) );
  OAI22_X1 U50 ( .A1(n83), .A2(n36), .B1(n43), .B2(n55), .ZN(n18) );
  INV_X1 U51 ( .A(D[14]), .ZN(n55) );
  OAI22_X1 U52 ( .A1(n80), .A2(n36), .B1(n44), .B2(n60), .ZN(n15) );
  INV_X1 U53 ( .A(D[17]), .ZN(n60) );
  OAI22_X1 U54 ( .A1(n76), .A2(n36), .B1(n45), .B2(n64), .ZN(n11) );
  INV_X1 U55 ( .A(D[21]), .ZN(n64) );
  OAI22_X1 U56 ( .A1(n90), .A2(n37), .B1(n41), .B2(n106), .ZN(n25) );
  INV_X1 U57 ( .A(D[7]), .ZN(n106) );
  OAI22_X1 U58 ( .A1(n94), .A2(n37), .B1(n40), .B2(n110), .ZN(n29) );
  INV_X1 U59 ( .A(D[3]), .ZN(n110) );
  OAI22_X1 U60 ( .A1(n97), .A2(n37), .B1(n39), .B2(n113), .ZN(n32) );
  INV_X1 U61 ( .A(D[0]), .ZN(n113) );
  OAI22_X1 U62 ( .A1(n96), .A2(n36), .B1(n39), .B2(n112), .ZN(n31) );
  INV_X1 U63 ( .A(D[1]), .ZN(n112) );
  OAI22_X1 U64 ( .A1(n95), .A2(n37), .B1(n40), .B2(n111), .ZN(n30) );
  INV_X1 U65 ( .A(D[2]), .ZN(n111) );
  OAI22_X1 U66 ( .A1(n93), .A2(n37), .B1(n40), .B2(n109), .ZN(n28) );
  INV_X1 U67 ( .A(D[4]), .ZN(n109) );
  OAI22_X1 U68 ( .A1(n92), .A2(n37), .B1(n41), .B2(n108), .ZN(n27) );
  INV_X1 U69 ( .A(D[5]), .ZN(n108) );
  OAI22_X1 U70 ( .A1(n91), .A2(n37), .B1(n41), .B2(n107), .ZN(n26) );
  INV_X1 U71 ( .A(D[6]), .ZN(n107) );
  OAI22_X1 U72 ( .A1(n89), .A2(n37), .B1(n41), .B2(n53), .ZN(n24) );
  INV_X1 U73 ( .A(D[8]), .ZN(n53) );
  OAI22_X1 U74 ( .A1(n87), .A2(n37), .B1(n42), .B2(n51), .ZN(n22) );
  INV_X1 U75 ( .A(D[10]), .ZN(n51) );
  OAI22_X1 U76 ( .A1(n86), .A2(n37), .B1(n42), .B2(n50), .ZN(n21) );
  INV_X1 U77 ( .A(D[11]), .ZN(n50) );
  OAI22_X1 U78 ( .A1(n88), .A2(n37), .B1(n42), .B2(n52), .ZN(n23) );
  INV_X1 U79 ( .A(D[9]), .ZN(n52) );
  BUF_X1 U80 ( .A(Enable_n), .Z(n35) );
  BUF_X1 U81 ( .A(Enable_n), .Z(n33) );
  BUF_X1 U82 ( .A(Enable_n), .Z(n34) );
endmodule


module PG_block_0 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_0 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n2;

  AOI21_X1 U1 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(G_out) );
endmodule


module PG_block_127 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_126 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_125 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_124 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_123 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_122 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_121 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_120 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_119 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_118 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_117 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_116 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_115 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_114 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_113 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_112 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_111 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_110 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_109 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_108 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_107 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_106 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_105 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_104 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_103 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_102 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_101 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_100 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_99 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_98 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_97 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_39 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_0 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n2;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n2), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n2) );
endmodule


module GENERAL_G_38 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_107 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_106 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_105 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_104 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_103 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_102 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_101 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_100 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_99 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_98 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_97 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_96 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_95 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_94 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_93 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_92 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_91 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_90 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_89 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_88 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_87 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_G_37 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_86 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_36 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_35 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_85 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_84 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_83 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_82 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_34 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_33 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_32 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_31 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   Cin, first_generate, \p_vett[4][3] , \p_vett[4][2] , \p_vett[3][3] ,
         \p_vett[3][2] , \p_vett[3][1] , \p_vett[2][7] , \p_vett[2][6] ,
         \p_vett[2][5] , \p_vett[2][4] , \p_vett[2][3] , \p_vett[2][2] ,
         \p_vett[2][1] , \p_vett[1][15] , \p_vett[1][14] , \p_vett[1][13] ,
         \p_vett[1][12] , \p_vett[1][11] , \p_vett[1][10] , \p_vett[1][9] ,
         \p_vett[1][8] , \p_vett[1][7] , \p_vett[1][6] , \p_vett[1][5] ,
         \p_vett[1][4] , \p_vett[1][3] , \p_vett[1][2] , \p_vett[1][1] ,
         \p_vett[0][31] , \p_vett[0][30] , \p_vett[0][29] , \p_vett[0][28] ,
         \p_vett[0][27] , \p_vett[0][26] , \p_vett[0][25] , \p_vett[0][24] ,
         \p_vett[0][23] , \p_vett[0][22] , \p_vett[0][21] , \p_vett[0][20] ,
         \p_vett[0][19] , \p_vett[0][18] , \p_vett[0][17] , \p_vett[0][16] ,
         \p_vett[0][15] , \p_vett[0][14] , \p_vett[0][13] , \p_vett[0][12] ,
         \p_vett[0][11] , \p_vett[0][10] , \p_vett[0][9] , \p_vett[0][8] ,
         \p_vett[0][7] , \p_vett[0][6] , \p_vett[0][5] , \p_vett[0][4] ,
         \p_vett[0][3] , \p_vett[0][2] , \p_vett[0][1] , \p_vett[0][0] ,
         \g_vett[4][3] , \g_vett[4][2] , \g_vett[3][3] , \g_vett[3][2] ,
         \g_vett[3][1] , \g_vett[2][7] , \g_vett[2][6] , \g_vett[2][5] ,
         \g_vett[2][4] , \g_vett[2][3] , \g_vett[2][2] , \g_vett[2][1] ,
         \g_vett[1][15] , \g_vett[1][14] , \g_vett[1][13] , \g_vett[1][12] ,
         \g_vett[1][11] , \g_vett[1][10] , \g_vett[1][9] , \g_vett[1][8] ,
         \g_vett[1][7] , \g_vett[1][6] , \g_vett[1][5] , \g_vett[1][4] ,
         \g_vett[1][3] , \g_vett[1][2] , \g_vett[1][1] , \g_vett[1][0] ,
         \g_vett[0][31] , \g_vett[0][30] , \g_vett[0][29] , \g_vett[0][28] ,
         \g_vett[0][27] , \g_vett[0][26] , \g_vett[0][25] , \g_vett[0][24] ,
         \g_vett[0][23] , \g_vett[0][22] , \g_vett[0][21] , \g_vett[0][20] ,
         \g_vett[0][19] , \g_vett[0][18] , \g_vett[0][17] , \g_vett[0][16] ,
         \g_vett[0][15] , \g_vett[0][14] , \g_vett[0][13] , \g_vett[0][12] ,
         \g_vett[0][11] , \g_vett[0][10] , \g_vett[0][9] , \g_vett[0][8] ,
         \g_vett[0][7] , \g_vett[0][6] , \g_vett[0][5] , \g_vett[0][4] ,
         \g_vett[0][3] , \g_vett[0][2] , \g_vett[0][1] , \g_vett[0][0] ;
  assign Co[0] = Cin;

  PG_block_0 PGblock_first ( .A(A[0]), .B(B[0]), .G(first_generate), .P(
        \p_vett[0][0] ) );
  GENERAL_G_0 G_first ( .G_in(first_generate), .P_in(\p_vett[0][0] ), 
        .G_in_prev(Cin), .G_out(\g_vett[0][0] ) );
  PG_block_127 PG_0_1 ( .A(A[1]), .B(B[1]), .G(\g_vett[0][1] ), .P(
        \p_vett[0][1] ) );
  PG_block_126 PG_0_2 ( .A(A[2]), .B(B[2]), .G(\g_vett[0][2] ), .P(
        \p_vett[0][2] ) );
  PG_block_125 PG_0_3 ( .A(A[3]), .B(B[3]), .G(\g_vett[0][3] ), .P(
        \p_vett[0][3] ) );
  PG_block_124 PG_0_4 ( .A(A[4]), .B(B[4]), .G(\g_vett[0][4] ), .P(
        \p_vett[0][4] ) );
  PG_block_123 PG_0_5 ( .A(A[5]), .B(B[5]), .G(\g_vett[0][5] ), .P(
        \p_vett[0][5] ) );
  PG_block_122 PG_0_6 ( .A(A[6]), .B(B[6]), .G(\g_vett[0][6] ), .P(
        \p_vett[0][6] ) );
  PG_block_121 PG_0_7 ( .A(A[7]), .B(B[7]), .G(\g_vett[0][7] ), .P(
        \p_vett[0][7] ) );
  PG_block_120 PG_0_8 ( .A(A[8]), .B(B[8]), .G(\g_vett[0][8] ), .P(
        \p_vett[0][8] ) );
  PG_block_119 PG_0_9 ( .A(A[9]), .B(B[9]), .G(\g_vett[0][9] ), .P(
        \p_vett[0][9] ) );
  PG_block_118 PG_0_10 ( .A(A[10]), .B(B[10]), .G(\g_vett[0][10] ), .P(
        \p_vett[0][10] ) );
  PG_block_117 PG_0_11 ( .A(A[11]), .B(B[11]), .G(\g_vett[0][11] ), .P(
        \p_vett[0][11] ) );
  PG_block_116 PG_0_12 ( .A(A[12]), .B(B[12]), .G(\g_vett[0][12] ), .P(
        \p_vett[0][12] ) );
  PG_block_115 PG_0_13 ( .A(A[13]), .B(B[13]), .G(\g_vett[0][13] ), .P(
        \p_vett[0][13] ) );
  PG_block_114 PG_0_14 ( .A(A[14]), .B(B[14]), .G(\g_vett[0][14] ), .P(
        \p_vett[0][14] ) );
  PG_block_113 PG_0_15 ( .A(A[15]), .B(B[15]), .G(\g_vett[0][15] ), .P(
        \p_vett[0][15] ) );
  PG_block_112 PG_0_16 ( .A(A[16]), .B(B[16]), .G(\g_vett[0][16] ), .P(
        \p_vett[0][16] ) );
  PG_block_111 PG_0_17 ( .A(A[17]), .B(B[17]), .G(\g_vett[0][17] ), .P(
        \p_vett[0][17] ) );
  PG_block_110 PG_0_18 ( .A(A[18]), .B(B[18]), .G(\g_vett[0][18] ), .P(
        \p_vett[0][18] ) );
  PG_block_109 PG_0_19 ( .A(A[19]), .B(B[19]), .G(\g_vett[0][19] ), .P(
        \p_vett[0][19] ) );
  PG_block_108 PG_0_20 ( .A(A[20]), .B(B[20]), .G(\g_vett[0][20] ), .P(
        \p_vett[0][20] ) );
  PG_block_107 PG_0_21 ( .A(A[21]), .B(B[21]), .G(\g_vett[0][21] ), .P(
        \p_vett[0][21] ) );
  PG_block_106 PG_0_22 ( .A(A[22]), .B(B[22]), .G(\g_vett[0][22] ), .P(
        \p_vett[0][22] ) );
  PG_block_105 PG_0_23 ( .A(A[23]), .B(B[23]), .G(\g_vett[0][23] ), .P(
        \p_vett[0][23] ) );
  PG_block_104 PG_0_24 ( .A(A[24]), .B(B[24]), .G(\g_vett[0][24] ), .P(
        \p_vett[0][24] ) );
  PG_block_103 PG_0_25 ( .A(A[25]), .B(B[25]), .G(\g_vett[0][25] ), .P(
        \p_vett[0][25] ) );
  PG_block_102 PG_0_26 ( .A(A[26]), .B(B[26]), .G(\g_vett[0][26] ), .P(
        \p_vett[0][26] ) );
  PG_block_101 PG_0_27 ( .A(A[27]), .B(B[27]), .G(\g_vett[0][27] ), .P(
        \p_vett[0][27] ) );
  PG_block_100 PG_0_28 ( .A(A[28]), .B(B[28]), .G(\g_vett[0][28] ), .P(
        \p_vett[0][28] ) );
  PG_block_99 PG_0_29 ( .A(A[29]), .B(B[29]), .G(\g_vett[0][29] ), .P(
        \p_vett[0][29] ) );
  PG_block_98 PG_0_30 ( .A(A[30]), .B(B[30]), .G(\g_vett[0][30] ), .P(
        \p_vett[0][30] ) );
  PG_block_97 PG_0_31 ( .A(A[31]), .B(B[31]), .G(\g_vett[0][31] ), .P(
        \p_vett[0][31] ) );
  GENERAL_G_39 G_0_0_0 ( .G_in(\g_vett[0][1] ), .P_in(\p_vett[0][1] ), 
        .G_in_prev(\g_vett[0][0] ), .G_out(\g_vett[1][0] ) );
  GENERAL_PG_0 PG_1_0_0 ( .G_in(\g_vett[0][3] ), .P_in(\p_vett[0][3] ), 
        .G_in_prev(\g_vett[0][2] ), .P_in_prev(\p_vett[0][2] ), .G_out(
        \g_vett[1][1] ), .P_out(\p_vett[1][1] ) );
  GENERAL_G_38 G_1_0_0 ( .G_in(\g_vett[1][1] ), .P_in(\p_vett[1][1] ), 
        .G_in_prev(\g_vett[1][0] ), .G_out(Co[1]) );
  GENERAL_PG_107 PG_2_0_1 ( .G_in(\g_vett[0][5] ), .P_in(\p_vett[0][5] ), 
        .G_in_prev(\g_vett[0][4] ), .P_in_prev(\p_vett[0][4] ), .G_out(
        \g_vett[1][2] ), .P_out(\p_vett[1][2] ) );
  GENERAL_PG_106 PG_3_0_1 ( .G_in(\g_vett[0][7] ), .P_in(\p_vett[0][7] ), 
        .G_in_prev(\g_vett[0][6] ), .P_in_prev(\p_vett[0][6] ), .G_out(
        \g_vett[1][3] ), .P_out(\p_vett[1][3] ) );
  GENERAL_PG_105 PG_4_0_1 ( .G_in(\g_vett[1][3] ), .P_in(\p_vett[1][3] ), 
        .G_in_prev(\g_vett[1][2] ), .P_in_prev(\p_vett[1][2] ), .G_out(
        \g_vett[2][1] ), .P_out(\p_vett[2][1] ) );
  GENERAL_PG_104 PG_2_0_2 ( .G_in(\g_vett[0][9] ), .P_in(\p_vett[0][9] ), 
        .G_in_prev(\g_vett[0][8] ), .P_in_prev(\p_vett[0][8] ), .G_out(
        \g_vett[1][4] ), .P_out(\p_vett[1][4] ) );
  GENERAL_PG_103 PG_3_0_2 ( .G_in(\g_vett[0][11] ), .P_in(\p_vett[0][11] ), 
        .G_in_prev(\g_vett[0][10] ), .P_in_prev(\p_vett[0][10] ), .G_out(
        \g_vett[1][5] ), .P_out(\p_vett[1][5] ) );
  GENERAL_PG_102 PG_4_0_2 ( .G_in(\g_vett[1][5] ), .P_in(\p_vett[1][5] ), 
        .G_in_prev(\g_vett[1][4] ), .P_in_prev(\p_vett[1][4] ), .G_out(
        \g_vett[2][2] ), .P_out(\p_vett[2][2] ) );
  GENERAL_PG_101 PG_2_0_3 ( .G_in(\g_vett[0][13] ), .P_in(\p_vett[0][13] ), 
        .G_in_prev(\g_vett[0][12] ), .P_in_prev(\p_vett[0][12] ), .G_out(
        \g_vett[1][6] ), .P_out(\p_vett[1][6] ) );
  GENERAL_PG_100 PG_3_0_3 ( .G_in(\g_vett[0][15] ), .P_in(\p_vett[0][15] ), 
        .G_in_prev(\g_vett[0][14] ), .P_in_prev(\p_vett[0][14] ), .G_out(
        \g_vett[1][7] ), .P_out(\p_vett[1][7] ) );
  GENERAL_PG_99 PG_4_0_3 ( .G_in(\g_vett[1][7] ), .P_in(\p_vett[1][7] ), 
        .G_in_prev(\g_vett[1][6] ), .P_in_prev(\p_vett[1][6] ), .G_out(
        \g_vett[2][3] ), .P_out(\p_vett[2][3] ) );
  GENERAL_PG_98 PG_2_0_4 ( .G_in(\g_vett[0][17] ), .P_in(\p_vett[0][17] ), 
        .G_in_prev(\g_vett[0][16] ), .P_in_prev(\p_vett[0][16] ), .G_out(
        \g_vett[1][8] ), .P_out(\p_vett[1][8] ) );
  GENERAL_PG_97 PG_3_0_4 ( .G_in(\g_vett[0][19] ), .P_in(\p_vett[0][19] ), 
        .G_in_prev(\g_vett[0][18] ), .P_in_prev(\p_vett[0][18] ), .G_out(
        \g_vett[1][9] ), .P_out(\p_vett[1][9] ) );
  GENERAL_PG_96 PG_4_0_4 ( .G_in(\g_vett[1][9] ), .P_in(\p_vett[1][9] ), 
        .G_in_prev(\g_vett[1][8] ), .P_in_prev(\p_vett[1][8] ), .G_out(
        \g_vett[2][4] ), .P_out(\p_vett[2][4] ) );
  GENERAL_PG_95 PG_2_0_5 ( .G_in(\g_vett[0][21] ), .P_in(\p_vett[0][21] ), 
        .G_in_prev(\g_vett[0][20] ), .P_in_prev(\p_vett[0][20] ), .G_out(
        \g_vett[1][10] ), .P_out(\p_vett[1][10] ) );
  GENERAL_PG_94 PG_3_0_5 ( .G_in(\g_vett[0][23] ), .P_in(\p_vett[0][23] ), 
        .G_in_prev(\g_vett[0][22] ), .P_in_prev(\p_vett[0][22] ), .G_out(
        \g_vett[1][11] ), .P_out(\p_vett[1][11] ) );
  GENERAL_PG_93 PG_4_0_5 ( .G_in(\g_vett[1][11] ), .P_in(\p_vett[1][11] ), 
        .G_in_prev(\g_vett[1][10] ), .P_in_prev(\p_vett[1][10] ), .G_out(
        \g_vett[2][5] ), .P_out(\p_vett[2][5] ) );
  GENERAL_PG_92 PG_2_0_6 ( .G_in(\g_vett[0][25] ), .P_in(\p_vett[0][25] ), 
        .G_in_prev(\g_vett[0][24] ), .P_in_prev(\p_vett[0][24] ), .G_out(
        \g_vett[1][12] ), .P_out(\p_vett[1][12] ) );
  GENERAL_PG_91 PG_3_0_6 ( .G_in(\g_vett[0][27] ), .P_in(\p_vett[0][27] ), 
        .G_in_prev(\g_vett[0][26] ), .P_in_prev(\p_vett[0][26] ), .G_out(
        \g_vett[1][13] ), .P_out(\p_vett[1][13] ) );
  GENERAL_PG_90 PG_4_0_6 ( .G_in(\g_vett[1][13] ), .P_in(\p_vett[1][13] ), 
        .G_in_prev(\g_vett[1][12] ), .P_in_prev(\p_vett[1][12] ), .G_out(
        \g_vett[2][6] ), .P_out(\p_vett[2][6] ) );
  GENERAL_PG_89 PG_2_0_7 ( .G_in(\g_vett[0][29] ), .P_in(\p_vett[0][29] ), 
        .G_in_prev(\g_vett[0][28] ), .P_in_prev(\p_vett[0][28] ), .G_out(
        \g_vett[1][14] ), .P_out(\p_vett[1][14] ) );
  GENERAL_PG_88 PG_3_0_7 ( .G_in(\g_vett[0][31] ), .P_in(\p_vett[0][31] ), 
        .G_in_prev(\g_vett[0][30] ), .P_in_prev(\p_vett[0][30] ), .G_out(
        \g_vett[1][15] ), .P_out(\p_vett[1][15] ) );
  GENERAL_PG_87 PG_4_0_7 ( .G_in(\g_vett[1][15] ), .P_in(\p_vett[1][15] ), 
        .G_in_prev(\g_vett[1][14] ), .P_in_prev(\p_vett[1][14] ), .G_out(
        \g_vett[2][7] ), .P_out(\p_vett[2][7] ) );
  GENERAL_G_37 G_2_1_0 ( .G_in(\g_vett[2][1] ), .P_in(\p_vett[2][1] ), 
        .G_in_prev(Co[1]), .G_out(Co[2]) );
  GENERAL_PG_86 PG_5_1_0 ( .G_in(\g_vett[2][3] ), .P_in(\p_vett[2][3] ), 
        .G_in_prev(\g_vett[2][2] ), .P_in_prev(\p_vett[2][2] ), .G_out(
        \g_vett[3][1] ), .P_out(\p_vett[3][1] ) );
  GENERAL_G_36 G_3_1_0 ( .G_in(\g_vett[2][2] ), .P_in(\p_vett[2][2] ), 
        .G_in_prev(Co[2]), .G_out(Co[3]) );
  GENERAL_G_35 G_4_1_0 ( .G_in(\g_vett[3][1] ), .P_in(\p_vett[3][1] ), 
        .G_in_prev(Co[2]), .G_out(Co[4]) );
  GENERAL_PG_85 PG_6_1_1 ( .G_in(\g_vett[2][5] ), .P_in(\p_vett[2][5] ), 
        .G_in_prev(\g_vett[2][4] ), .P_in_prev(\p_vett[2][4] ), .G_out(
        \g_vett[3][2] ), .P_out(\p_vett[3][2] ) );
  GENERAL_PG_84 PG_7_1_1 ( .G_in(\g_vett[2][7] ), .P_in(\p_vett[2][7] ), 
        .G_in_prev(\g_vett[2][6] ), .P_in_prev(\p_vett[2][6] ), .G_out(
        \g_vett[3][3] ), .P_out(\p_vett[3][3] ) );
  GENERAL_PG_83 PG_8_1_1 ( .G_in(\g_vett[2][6] ), .P_in(\p_vett[2][6] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][2] ), .P_out(\p_vett[4][2] ) );
  GENERAL_PG_82 PG_9_1_1 ( .G_in(\g_vett[3][3] ), .P_in(\p_vett[3][3] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][3] ), .P_out(\p_vett[4][3] ) );
  GENERAL_G_34 G_5_2_0 ( .G_in(\g_vett[2][4] ), .P_in(\p_vett[2][4] ), 
        .G_in_prev(Co[4]), .G_out(Co[5]) );
  GENERAL_G_33 G_6_2_1 ( .G_in(\g_vett[3][2] ), .P_in(\p_vett[3][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[6]) );
  GENERAL_G_32 G_7_2_2 ( .G_in(\g_vett[4][2] ), .P_in(\p_vett[4][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[7]) );
  GENERAL_G_31 G_8_2_3 ( .G_in(\g_vett[4][3] ), .P_in(\p_vett[4][3] ), 
        .G_in_prev(Co[4]) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n2) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_255 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_254 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_253 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_63 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_252 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_251 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_250 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_249 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n13;

  INV_X1 U1 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n9) );
  INV_X1 U3 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n8) );
  INV_X1 U5 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n7) );
  INV_X1 U7 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n6) );
  INV_X1 U9 ( .A(SEL), .ZN(n13) );
endmodule


module MUX21_GENERIC_NBIT4_63 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n13;

  INV_X1 U1 ( .A(n9), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n8), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n7), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n9) );
  INV_X1 U6 ( .A(SEL), .ZN(n13) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n8) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n7) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n6) );
endmodule


module CSblock_NBIT4_0 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_0 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_63 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_0 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_63 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_62 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_248 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_247 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_246 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_245 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_61 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_244 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_243 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_242 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_241 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_62 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_61 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_31 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_62 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_61 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_62 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_61 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_60 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_240 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_239 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_238 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_237 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_59 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_236 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_235 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_234 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_233 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_60 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_59 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_30 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_60 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_59 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_60 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_59 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_58 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_232 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_231 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_230 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_229 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_57 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_228 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_227 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_226 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_225 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_58 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_57 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_29 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_58 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_57 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_58 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_57 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_56 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_224 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_223 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_222 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_221 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_55 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_220 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_219 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_218 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_217 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_56 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U6 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_55 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_28 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_56 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_55 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_56 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_55 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_54 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_216 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_215 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_214 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_213 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_53 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_212 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_211 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_210 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_209 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_54 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_53 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_27 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_54 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_53 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_54 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_53 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_52 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_208 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_207 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_206 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_205 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_51 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_204 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_203 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_202 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_201 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_52 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_51 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_26 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_52 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_51 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_52 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_51 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_50 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_200 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_199 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_198 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_197 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_49 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_196 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_195 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_194 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_193 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_50 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_49 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_25 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_50 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_49 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_50 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_49 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module SUMGEN_NBIT32_NBLOCKS8_0 ( A, B, cin_vect, Co, SUM );
  input [31:0] A;
  input [31:0] B;
  input [7:0] cin_vect;
  output [31:0] SUM;
  output Co;


  CSblock_NBIT4_0 block_i_0 ( .A(A[3:0]), .B(B[3:0]), .cin(cin_vect[0]), .Y(
        SUM[3:0]) );
  CSblock_NBIT4_31 block_i_1 ( .A(A[7:4]), .B(B[7:4]), .cin(cin_vect[1]), .Y(
        SUM[7:4]) );
  CSblock_NBIT4_30 block_i_2 ( .A(A[11:8]), .B(B[11:8]), .cin(cin_vect[2]), 
        .Y(SUM[11:8]) );
  CSblock_NBIT4_29 block_i_3 ( .A(A[15:12]), .B(B[15:12]), .cin(cin_vect[3]), 
        .Y(SUM[15:12]) );
  CSblock_NBIT4_28 block_i_4 ( .A(A[19:16]), .B(B[19:16]), .cin(cin_vect[4]), 
        .Y(SUM[19:16]) );
  CSblock_NBIT4_27 block_i_5 ( .A(A[23:20]), .B(B[23:20]), .cin(cin_vect[5]), 
        .Y(SUM[23:20]) );
  CSblock_NBIT4_26 block_i_6 ( .A(A[27:24]), .B(B[27:24]), .cin(cin_vect[6]), 
        .Y(SUM[27:24]) );
  CSblock_NBIT4_25 block_i_7 ( .A(A[31:28]), .B(B[31:28]), .cin(cin_vect[7]), 
        .Y(SUM[31:28]), .Co(Co) );
endmodule


module P4_ADDER_NBIT32_NBIT_PER_BLOCK4_0 ( A, B, Cin, Cout, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input Cin;
  output Cout;

  wire   [7:0] outCarryGen;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 CG ( .A(A), .B(B), .Cin(Cin), .Co(
        outCarryGen) );
  SUMGEN_NBIT32_NBLOCKS8_0 SG ( .A(A), .B(B), .cin_vect(outCarryGen), .Co(Cout), .SUM(Y) );
endmodule


module REG_GEN_NBIT32_18 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n47), .Q(Q[31]), .QN(n145) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n47), .Q(Q[30]), .QN(n144) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n47), .Q(Q[29]), .QN(n143) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n47), .Q(Q[28]), .QN(n142) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n47), .Q(Q[27]), .QN(n141) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n47), .Q(Q[26]), .QN(n140) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n47), .Q(Q[25]), .QN(n139) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n47), .Q(Q[24]), .QN(n138) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n47), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n47), .Q(Q[22]), .QN(n136) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n47), .Q(Q[21]), .QN(n135) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n47), .Q(Q[20]), .QN(n134) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n48), .Q(Q[19]), .QN(n133) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n48), .Q(Q[18]), .QN(n132) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n48), .Q(Q[17]), .QN(n131) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n48), .Q(Q[16]), .QN(n130) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n48), .Q(Q[15]), .QN(n129) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n48), .Q(Q[14]), .QN(n128) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n48), .Q(Q[13]), .QN(n127) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n48), .Q(Q[12]), .QN(n126) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n48), .Q(Q[11]), .QN(n125) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n48), .Q(Q[10]), .QN(n124) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n48), .Q(Q[9]), .QN(n123) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n48), .Q(Q[8]), .QN(n122) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n49), .Q(Q[7]), .QN(n121) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n49), .Q(Q[6]), .QN(n120) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n49), .Q(Q[5]), .QN(n119) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n49), .Q(Q[4]), .QN(n118) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n49), .Q(Q[3]), .QN(n117) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n49), .Q(Q[2]), .QN(n116) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n49), .Q(Q[1]), .QN(n115) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n49), .Q(Q[0]), .QN(n114) );
  BUF_X1 U2 ( .A(RESET_n), .Z(n48) );
  BUF_X1 U3 ( .A(RESET_n), .Z(n47) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n49) );
  INV_X1 U5 ( .A(n46), .ZN(n37) );
  INV_X1 U6 ( .A(n46), .ZN(n36) );
  BUF_X1 U7 ( .A(n35), .Z(n46) );
  BUF_X1 U8 ( .A(n34), .Z(n41) );
  BUF_X1 U9 ( .A(n34), .Z(n42) );
  BUF_X1 U10 ( .A(n35), .Z(n44) );
  BUF_X1 U11 ( .A(n33), .Z(n38) );
  BUF_X1 U12 ( .A(n33), .Z(n39) );
  BUF_X1 U13 ( .A(n33), .Z(n40) );
  BUF_X1 U14 ( .A(n34), .Z(n43) );
  BUF_X1 U15 ( .A(n35), .Z(n45) );
  OAI22_X1 U16 ( .A1(n114), .A2(n37), .B1(n39), .B2(n113), .ZN(n32) );
  INV_X1 U17 ( .A(D[0]), .ZN(n113) );
  OAI22_X1 U18 ( .A1(n115), .A2(n36), .B1(n39), .B2(n112), .ZN(n31) );
  INV_X1 U19 ( .A(D[1]), .ZN(n112) );
  OAI22_X1 U20 ( .A1(n116), .A2(n37), .B1(n40), .B2(n111), .ZN(n30) );
  INV_X1 U21 ( .A(D[2]), .ZN(n111) );
  OAI22_X1 U22 ( .A1(n117), .A2(n37), .B1(n40), .B2(n110), .ZN(n29) );
  INV_X1 U23 ( .A(D[3]), .ZN(n110) );
  OAI22_X1 U24 ( .A1(n134), .A2(n36), .B1(n45), .B2(n65), .ZN(n12) );
  INV_X1 U25 ( .A(D[20]), .ZN(n65) );
  OAI22_X1 U26 ( .A1(n135), .A2(n36), .B1(n45), .B2(n64), .ZN(n11) );
  INV_X1 U27 ( .A(D[21]), .ZN(n64) );
  OAI22_X1 U28 ( .A1(n136), .A2(n36), .B1(n45), .B2(n63), .ZN(n10) );
  INV_X1 U29 ( .A(D[22]), .ZN(n63) );
  OAI22_X1 U30 ( .A1(n137), .A2(n37), .B1(n38), .B2(n62), .ZN(n9) );
  INV_X1 U31 ( .A(D[23]), .ZN(n62) );
  OAI22_X1 U32 ( .A1(n138), .A2(n37), .B1(n38), .B2(n101), .ZN(n8) );
  INV_X1 U33 ( .A(D[24]), .ZN(n101) );
  OAI22_X1 U34 ( .A1(n139), .A2(n36), .B1(n38), .B2(n100), .ZN(n7) );
  INV_X1 U35 ( .A(D[25]), .ZN(n100) );
  OAI22_X1 U36 ( .A1(n140), .A2(n37), .B1(n38), .B2(n99), .ZN(n6) );
  INV_X1 U37 ( .A(D[26]), .ZN(n99) );
  OAI22_X1 U38 ( .A1(n141), .A2(n36), .B1(n39), .B2(n98), .ZN(n5) );
  INV_X1 U39 ( .A(D[27]), .ZN(n98) );
  OAI22_X1 U40 ( .A1(n142), .A2(n36), .B1(n39), .B2(n105), .ZN(n4) );
  INV_X1 U41 ( .A(D[28]), .ZN(n105) );
  OAI22_X1 U42 ( .A1(n143), .A2(n37), .B1(n40), .B2(n104), .ZN(n3) );
  INV_X1 U43 ( .A(D[29]), .ZN(n104) );
  OAI22_X1 U44 ( .A1(n144), .A2(n36), .B1(n43), .B2(n103), .ZN(n2) );
  INV_X1 U45 ( .A(D[30]), .ZN(n103) );
  OAI22_X1 U46 ( .A1(n145), .A2(n36), .B1(n45), .B2(n102), .ZN(n1) );
  INV_X1 U47 ( .A(D[31]), .ZN(n102) );
  OAI22_X1 U48 ( .A1(n130), .A2(n36), .B1(n44), .B2(n61), .ZN(n16) );
  INV_X1 U49 ( .A(D[16]), .ZN(n61) );
  OAI22_X1 U50 ( .A1(n131), .A2(n36), .B1(n44), .B2(n60), .ZN(n15) );
  INV_X1 U51 ( .A(D[17]), .ZN(n60) );
  OAI22_X1 U52 ( .A1(n132), .A2(n36), .B1(n44), .B2(n59), .ZN(n14) );
  INV_X1 U53 ( .A(D[18]), .ZN(n59) );
  OAI22_X1 U54 ( .A1(n122), .A2(n37), .B1(n41), .B2(n53), .ZN(n24) );
  INV_X1 U55 ( .A(D[8]), .ZN(n53) );
  OAI22_X1 U56 ( .A1(n123), .A2(n37), .B1(n42), .B2(n52), .ZN(n23) );
  INV_X1 U57 ( .A(D[9]), .ZN(n52) );
  OAI22_X1 U58 ( .A1(n124), .A2(n37), .B1(n42), .B2(n51), .ZN(n22) );
  INV_X1 U59 ( .A(D[10]), .ZN(n51) );
  OAI22_X1 U60 ( .A1(n133), .A2(n36), .B1(n44), .B2(n58), .ZN(n13) );
  INV_X1 U61 ( .A(D[19]), .ZN(n58) );
  OAI22_X1 U62 ( .A1(n118), .A2(n37), .B1(n40), .B2(n109), .ZN(n28) );
  INV_X1 U63 ( .A(D[4]), .ZN(n109) );
  OAI22_X1 U64 ( .A1(n119), .A2(n37), .B1(n41), .B2(n108), .ZN(n27) );
  INV_X1 U65 ( .A(D[5]), .ZN(n108) );
  OAI22_X1 U66 ( .A1(n120), .A2(n37), .B1(n41), .B2(n107), .ZN(n26) );
  INV_X1 U67 ( .A(D[6]), .ZN(n107) );
  OAI22_X1 U68 ( .A1(n126), .A2(n37), .B1(n42), .B2(n57), .ZN(n20) );
  INV_X1 U69 ( .A(D[12]), .ZN(n57) );
  OAI22_X1 U70 ( .A1(n127), .A2(n36), .B1(n43), .B2(n56), .ZN(n19) );
  INV_X1 U71 ( .A(D[13]), .ZN(n56) );
  OAI22_X1 U72 ( .A1(n128), .A2(n36), .B1(n43), .B2(n55), .ZN(n18) );
  INV_X1 U73 ( .A(D[14]), .ZN(n55) );
  OAI22_X1 U74 ( .A1(n125), .A2(n37), .B1(n42), .B2(n50), .ZN(n21) );
  INV_X1 U75 ( .A(D[11]), .ZN(n50) );
  OAI22_X1 U76 ( .A1(n121), .A2(n37), .B1(n41), .B2(n106), .ZN(n25) );
  INV_X1 U77 ( .A(D[7]), .ZN(n106) );
  OAI22_X1 U78 ( .A1(n129), .A2(n36), .B1(n43), .B2(n54), .ZN(n17) );
  INV_X1 U79 ( .A(D[15]), .ZN(n54) );
  BUF_X1 U80 ( .A(Enable_n), .Z(n35) );
  BUF_X1 U81 ( .A(Enable_n), .Z(n33) );
  BUF_X1 U82 ( .A(Enable_n), .Z(n34) );
endmodule


module REG_GEN_NBIT32_17 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n49), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n49), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n49), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n49), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n49), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n49), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n49), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n49), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n48), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n48), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n48), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n48), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n48), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n48), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n48), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n48), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n48), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n48), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n48), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n48), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n47), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n47), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n47), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n47), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n47), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n47), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n47), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n47), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n47), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n47), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n47), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n47), .Q(Q[0]), .QN(n97) );
  BUF_X1 U2 ( .A(RESET_n), .Z(n47) );
  BUF_X1 U3 ( .A(RESET_n), .Z(n48) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n49) );
  INV_X1 U5 ( .A(n46), .ZN(n37) );
  INV_X1 U6 ( .A(n46), .ZN(n36) );
  BUF_X1 U7 ( .A(n35), .Z(n46) );
  BUF_X1 U8 ( .A(n34), .Z(n41) );
  BUF_X1 U9 ( .A(n34), .Z(n42) );
  BUF_X1 U10 ( .A(n35), .Z(n44) );
  BUF_X1 U11 ( .A(n33), .Z(n38) );
  BUF_X1 U12 ( .A(n33), .Z(n39) );
  BUF_X1 U13 ( .A(n33), .Z(n40) );
  BUF_X1 U14 ( .A(n34), .Z(n43) );
  BUF_X1 U15 ( .A(n35), .Z(n45) );
  OAI22_X1 U16 ( .A1(n97), .A2(n37), .B1(n39), .B2(n113), .ZN(n32) );
  INV_X1 U17 ( .A(D[0]), .ZN(n113) );
  OAI22_X1 U18 ( .A1(n96), .A2(n36), .B1(n39), .B2(n112), .ZN(n31) );
  INV_X1 U19 ( .A(D[1]), .ZN(n112) );
  OAI22_X1 U20 ( .A1(n95), .A2(n37), .B1(n40), .B2(n111), .ZN(n30) );
  INV_X1 U21 ( .A(D[2]), .ZN(n111) );
  OAI22_X1 U22 ( .A1(n94), .A2(n37), .B1(n40), .B2(n110), .ZN(n29) );
  INV_X1 U23 ( .A(D[3]), .ZN(n110) );
  OAI22_X1 U24 ( .A1(n93), .A2(n37), .B1(n40), .B2(n109), .ZN(n28) );
  INV_X1 U25 ( .A(D[4]), .ZN(n109) );
  OAI22_X1 U26 ( .A1(n92), .A2(n37), .B1(n41), .B2(n108), .ZN(n27) );
  INV_X1 U27 ( .A(D[5]), .ZN(n108) );
  OAI22_X1 U28 ( .A1(n91), .A2(n37), .B1(n41), .B2(n107), .ZN(n26) );
  INV_X1 U29 ( .A(D[6]), .ZN(n107) );
  OAI22_X1 U30 ( .A1(n90), .A2(n37), .B1(n41), .B2(n106), .ZN(n25) );
  INV_X1 U31 ( .A(D[7]), .ZN(n106) );
  OAI22_X1 U32 ( .A1(n89), .A2(n37), .B1(n41), .B2(n105), .ZN(n24) );
  INV_X1 U33 ( .A(D[8]), .ZN(n105) );
  OAI22_X1 U34 ( .A1(n88), .A2(n37), .B1(n42), .B2(n104), .ZN(n23) );
  INV_X1 U35 ( .A(D[9]), .ZN(n104) );
  OAI22_X1 U36 ( .A1(n87), .A2(n37), .B1(n42), .B2(n103), .ZN(n22) );
  INV_X1 U37 ( .A(D[10]), .ZN(n103) );
  OAI22_X1 U38 ( .A1(n86), .A2(n37), .B1(n42), .B2(n102), .ZN(n21) );
  INV_X1 U39 ( .A(D[11]), .ZN(n102) );
  OAI22_X1 U40 ( .A1(n85), .A2(n37), .B1(n42), .B2(n101), .ZN(n20) );
  INV_X1 U41 ( .A(D[12]), .ZN(n101) );
  OAI22_X1 U42 ( .A1(n84), .A2(n36), .B1(n43), .B2(n100), .ZN(n19) );
  INV_X1 U43 ( .A(D[13]), .ZN(n100) );
  OAI22_X1 U44 ( .A1(n83), .A2(n36), .B1(n43), .B2(n99), .ZN(n18) );
  INV_X1 U45 ( .A(D[14]), .ZN(n99) );
  OAI22_X1 U46 ( .A1(n82), .A2(n36), .B1(n43), .B2(n98), .ZN(n17) );
  INV_X1 U47 ( .A(D[15]), .ZN(n98) );
  OAI22_X1 U48 ( .A1(n81), .A2(n36), .B1(n44), .B2(n65), .ZN(n16) );
  INV_X1 U49 ( .A(D[16]), .ZN(n65) );
  OAI22_X1 U50 ( .A1(n80), .A2(n36), .B1(n44), .B2(n64), .ZN(n15) );
  INV_X1 U51 ( .A(D[17]), .ZN(n64) );
  OAI22_X1 U52 ( .A1(n79), .A2(n36), .B1(n44), .B2(n63), .ZN(n14) );
  INV_X1 U53 ( .A(D[18]), .ZN(n63) );
  OAI22_X1 U54 ( .A1(n78), .A2(n36), .B1(n44), .B2(n62), .ZN(n13) );
  INV_X1 U55 ( .A(D[19]), .ZN(n62) );
  OAI22_X1 U56 ( .A1(n77), .A2(n36), .B1(n45), .B2(n61), .ZN(n12) );
  INV_X1 U57 ( .A(D[20]), .ZN(n61) );
  OAI22_X1 U58 ( .A1(n76), .A2(n36), .B1(n45), .B2(n60), .ZN(n11) );
  INV_X1 U59 ( .A(D[21]), .ZN(n60) );
  OAI22_X1 U60 ( .A1(n75), .A2(n36), .B1(n45), .B2(n59), .ZN(n10) );
  INV_X1 U61 ( .A(D[22]), .ZN(n59) );
  OAI22_X1 U62 ( .A1(n74), .A2(n37), .B1(n38), .B2(n58), .ZN(n9) );
  INV_X1 U63 ( .A(D[23]), .ZN(n58) );
  OAI22_X1 U64 ( .A1(n73), .A2(n36), .B1(n38), .B2(n57), .ZN(n8) );
  INV_X1 U65 ( .A(D[24]), .ZN(n57) );
  OAI22_X1 U66 ( .A1(n72), .A2(n37), .B1(n38), .B2(n56), .ZN(n7) );
  INV_X1 U67 ( .A(D[25]), .ZN(n56) );
  OAI22_X1 U68 ( .A1(n71), .A2(n36), .B1(n38), .B2(n55), .ZN(n6) );
  INV_X1 U69 ( .A(D[26]), .ZN(n55) );
  OAI22_X1 U70 ( .A1(n70), .A2(n37), .B1(n39), .B2(n54), .ZN(n5) );
  INV_X1 U71 ( .A(D[27]), .ZN(n54) );
  OAI22_X1 U72 ( .A1(n69), .A2(n36), .B1(n39), .B2(n53), .ZN(n4) );
  INV_X1 U73 ( .A(D[28]), .ZN(n53) );
  OAI22_X1 U74 ( .A1(n68), .A2(n37), .B1(n40), .B2(n52), .ZN(n3) );
  INV_X1 U75 ( .A(D[29]), .ZN(n52) );
  OAI22_X1 U76 ( .A1(n67), .A2(n36), .B1(n43), .B2(n51), .ZN(n2) );
  INV_X1 U77 ( .A(D[30]), .ZN(n51) );
  OAI22_X1 U78 ( .A1(n66), .A2(n36), .B1(n45), .B2(n50), .ZN(n1) );
  INV_X1 U79 ( .A(D[31]), .ZN(n50) );
  BUF_X1 U80 ( .A(Enable_n), .Z(n35) );
  BUF_X1 U81 ( .A(Enable_n), .Z(n33) );
  BUF_X1 U82 ( .A(Enable_n), .Z(n34) );
endmodule


module fetchUnit_nbit32 ( Clk, Rst, en_reg, PC_branch_jump, dout_IRAM, PC_op, 
        PC_Next_out, addr_IRAM, IRAM_reg_out );
  input [31:0] PC_branch_jump;
  input [31:0] dout_IRAM;
  output [31:0] PC_Next_out;
  output [31:0] addr_IRAM;
  output [31:0] IRAM_reg_out;
  input Clk, Rst, en_reg, PC_op;

  wire   [31:0] PC_Next;
  wire   [31:0] PC_in;

  MUX21_GENERIC_NBIT32_0 mux_PC ( .A(PC_Next), .B(PC_branch_jump), .SEL(PC_op), 
        .Y(PC_in) );
  REG_GEN_NBIT32_0 PC_block ( .D(PC_in), .CK(Clk), .Enable_n(en_reg), 
        .RESET_n(Rst), .Q(addr_IRAM) );
  P4_ADDER_NBIT32_NBIT_PER_BLOCK4_0 PC_ADD ( .A(addr_IRAM), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .Cin(1'b0), .Y(PC_Next) );
  REG_GEN_NBIT32_18 IF_reg_PC_Next ( .D(PC_Next), .CK(Clk), .Enable_n(en_reg), 
        .RESET_n(Rst), .Q(PC_Next_out) );
  REG_GEN_NBIT32_17 IF_reg_IRAM_out ( .D(dout_IRAM), .CK(Clk), .Enable_n(
        en_reg), .RESET_n(Rst), .Q(IRAM_reg_out) );
endmodule


module sign_extension_sign_init26_sign_ext32 ( data_in, data_out );
  input [25:0] data_in;
  output [31:0] data_out;
  wire   data_out_31;
  assign data_out[31] = data_out_31;
  assign data_out[30] = data_out_31;
  assign data_out[29] = data_out_31;
  assign data_out[28] = data_out_31;
  assign data_out[27] = data_out_31;
  assign data_out[26] = data_out_31;
  assign data_out[25] = data_out_31;
  assign data_out_31 = data_in[25];
  assign data_out[24] = data_in[24];
  assign data_out[23] = data_in[23];
  assign data_out[22] = data_in[22];
  assign data_out[21] = data_in[21];
  assign data_out[20] = data_in[20];
  assign data_out[19] = data_in[19];
  assign data_out[18] = data_in[18];
  assign data_out[17] = data_in[17];
  assign data_out[16] = data_in[16];
  assign data_out[15] = data_in[15];
  assign data_out[14] = data_in[14];
  assign data_out[13] = data_in[13];
  assign data_out[12] = data_in[12];
  assign data_out[11] = data_in[11];
  assign data_out[10] = data_in[10];
  assign data_out[9] = data_in[9];
  assign data_out[8] = data_in[8];
  assign data_out[7] = data_in[7];
  assign data_out[6] = data_in[6];
  assign data_out[5] = data_in[5];
  assign data_out[4] = data_in[4];
  assign data_out[3] = data_in[3];
  assign data_out[2] = data_in[2];
  assign data_out[1] = data_in[1];
  assign data_out[0] = data_in[0];

endmodule


module register_file_nbit_reg32_n_reg32_nbit_addr5 ( reset, enable, rd1, rd2, 
        wr, add_wr, add_rd1, add_rd2, datain, out1, out2 );
  input [4:0] add_wr;
  input [4:0] add_rd1;
  input [4:0] add_rd2;
  input [31:0] datain;
  output [31:0] out1;
  output [31:0] out2;
  input reset, enable, rd1, rd2, wr;
  wire   \registers[1][31] , \registers[1][30] , \registers[1][29] ,
         \registers[1][28] , \registers[1][27] , \registers[1][26] ,
         \registers[1][25] , \registers[1][24] , \registers[1][23] ,
         \registers[1][22] , \registers[1][21] , \registers[1][20] ,
         \registers[1][19] , \registers[1][18] , \registers[1][17] ,
         \registers[1][16] , \registers[1][15] , \registers[1][14] ,
         \registers[1][13] , \registers[1][12] , \registers[1][11] ,
         \registers[1][10] , \registers[1][9] , \registers[1][8] ,
         \registers[1][7] , \registers[1][6] , \registers[1][5] ,
         \registers[1][4] , \registers[1][3] , \registers[1][2] ,
         \registers[1][1] , \registers[1][0] , \registers[2][31] ,
         \registers[2][30] , \registers[2][29] , \registers[2][28] ,
         \registers[2][27] , \registers[2][26] , \registers[2][25] ,
         \registers[2][24] , \registers[2][23] , \registers[2][22] ,
         \registers[2][21] , \registers[2][20] , \registers[2][19] ,
         \registers[2][18] , \registers[2][17] , \registers[2][16] ,
         \registers[2][15] , \registers[2][14] , \registers[2][13] ,
         \registers[2][12] , \registers[2][11] , \registers[2][10] ,
         \registers[2][9] , \registers[2][8] , \registers[2][7] ,
         \registers[2][6] , \registers[2][5] , \registers[2][4] ,
         \registers[2][3] , \registers[2][2] , \registers[2][1] ,
         \registers[2][0] , \registers[3][31] , \registers[3][30] ,
         \registers[3][29] , \registers[3][28] , \registers[3][27] ,
         \registers[3][26] , \registers[3][25] , \registers[3][24] ,
         \registers[3][23] , \registers[3][22] , \registers[3][21] ,
         \registers[3][20] , \registers[3][19] , \registers[3][18] ,
         \registers[3][17] , \registers[3][16] , \registers[3][15] ,
         \registers[3][14] , \registers[3][13] , \registers[3][12] ,
         \registers[3][11] , \registers[3][10] , \registers[3][9] ,
         \registers[3][8] , \registers[3][7] , \registers[3][6] ,
         \registers[3][5] , \registers[3][4] , \registers[3][3] ,
         \registers[3][2] , \registers[3][1] , \registers[3][0] ,
         \registers[4][31] , \registers[4][30] , \registers[4][29] ,
         \registers[4][28] , \registers[4][27] , \registers[4][26] ,
         \registers[4][25] , \registers[4][24] , \registers[4][23] ,
         \registers[4][22] , \registers[4][21] , \registers[4][20] ,
         \registers[4][19] , \registers[4][18] , \registers[4][17] ,
         \registers[4][16] , \registers[4][15] , \registers[4][14] ,
         \registers[4][13] , \registers[4][12] , \registers[4][11] ,
         \registers[4][10] , \registers[4][9] , \registers[4][8] ,
         \registers[4][7] , \registers[4][6] , \registers[4][5] ,
         \registers[4][4] , \registers[4][3] , \registers[4][2] ,
         \registers[4][1] , \registers[4][0] , \registers[5][31] ,
         \registers[5][30] , \registers[5][29] , \registers[5][28] ,
         \registers[5][27] , \registers[5][26] , \registers[5][25] ,
         \registers[5][24] , \registers[5][23] , \registers[5][22] ,
         \registers[5][21] , \registers[5][20] , \registers[5][19] ,
         \registers[5][18] , \registers[5][17] , \registers[5][16] ,
         \registers[5][15] , \registers[5][14] , \registers[5][13] ,
         \registers[5][12] , \registers[5][11] , \registers[5][10] ,
         \registers[5][9] , \registers[5][8] , \registers[5][7] ,
         \registers[5][6] , \registers[5][5] , \registers[5][4] ,
         \registers[5][3] , \registers[5][2] , \registers[5][1] ,
         \registers[5][0] , \registers[6][31] , \registers[6][30] ,
         \registers[6][29] , \registers[6][28] , \registers[6][27] ,
         \registers[6][26] , \registers[6][25] , \registers[6][24] ,
         \registers[6][23] , \registers[6][22] , \registers[6][21] ,
         \registers[6][20] , \registers[6][19] , \registers[6][18] ,
         \registers[6][17] , \registers[6][16] , \registers[6][15] ,
         \registers[6][14] , \registers[6][13] , \registers[6][12] ,
         \registers[6][11] , \registers[6][10] , \registers[6][9] ,
         \registers[6][8] , \registers[6][7] , \registers[6][6] ,
         \registers[6][5] , \registers[6][4] , \registers[6][3] ,
         \registers[6][2] , \registers[6][1] , \registers[6][0] ,
         \registers[7][31] , \registers[7][30] , \registers[7][29] ,
         \registers[7][28] , \registers[7][27] , \registers[7][26] ,
         \registers[7][25] , \registers[7][24] , \registers[7][23] ,
         \registers[7][22] , \registers[7][21] , \registers[7][20] ,
         \registers[7][19] , \registers[7][18] , \registers[7][17] ,
         \registers[7][16] , \registers[7][15] , \registers[7][14] ,
         \registers[7][13] , \registers[7][12] , \registers[7][11] ,
         \registers[7][10] , \registers[7][9] , \registers[7][8] ,
         \registers[7][7] , \registers[7][6] , \registers[7][5] ,
         \registers[7][4] , \registers[7][3] , \registers[7][2] ,
         \registers[7][1] , \registers[7][0] , \registers[8][31] ,
         \registers[8][30] , \registers[8][29] , \registers[8][28] ,
         \registers[8][27] , \registers[8][26] , \registers[8][25] ,
         \registers[8][24] , \registers[8][23] , \registers[8][22] ,
         \registers[8][21] , \registers[8][20] , \registers[8][19] ,
         \registers[8][18] , \registers[8][17] , \registers[8][16] ,
         \registers[8][15] , \registers[8][14] , \registers[8][13] ,
         \registers[8][12] , \registers[8][11] , \registers[8][10] ,
         \registers[8][9] , \registers[8][8] , \registers[8][7] ,
         \registers[8][6] , \registers[8][5] , \registers[8][4] ,
         \registers[8][3] , \registers[8][2] , \registers[8][1] ,
         \registers[8][0] , \registers[9][31] , \registers[9][30] ,
         \registers[9][29] , \registers[9][28] , \registers[9][27] ,
         \registers[9][26] , \registers[9][25] , \registers[9][24] ,
         \registers[9][23] , \registers[9][22] , \registers[9][21] ,
         \registers[9][20] , \registers[9][19] , \registers[9][18] ,
         \registers[9][17] , \registers[9][16] , \registers[9][15] ,
         \registers[9][14] , \registers[9][13] , \registers[9][12] ,
         \registers[9][11] , \registers[9][10] , \registers[9][9] ,
         \registers[9][8] , \registers[9][7] , \registers[9][6] ,
         \registers[9][5] , \registers[9][4] , \registers[9][3] ,
         \registers[9][2] , \registers[9][1] , \registers[9][0] ,
         \registers[10][31] , \registers[10][30] , \registers[10][29] ,
         \registers[10][28] , \registers[10][27] , \registers[10][26] ,
         \registers[10][25] , \registers[10][24] , \registers[10][23] ,
         \registers[10][22] , \registers[10][21] , \registers[10][20] ,
         \registers[10][19] , \registers[10][18] , \registers[10][17] ,
         \registers[10][16] , \registers[10][15] , \registers[10][14] ,
         \registers[10][13] , \registers[10][12] , \registers[10][11] ,
         \registers[10][10] , \registers[10][9] , \registers[10][8] ,
         \registers[10][7] , \registers[10][6] , \registers[10][5] ,
         \registers[10][4] , \registers[10][3] , \registers[10][2] ,
         \registers[10][1] , \registers[10][0] , \registers[11][31] ,
         \registers[11][30] , \registers[11][29] , \registers[11][28] ,
         \registers[11][27] , \registers[11][26] , \registers[11][25] ,
         \registers[11][24] , \registers[11][23] , \registers[11][22] ,
         \registers[11][21] , \registers[11][20] , \registers[11][19] ,
         \registers[11][18] , \registers[11][17] , \registers[11][16] ,
         \registers[11][15] , \registers[11][14] , \registers[11][13] ,
         \registers[11][12] , \registers[11][11] , \registers[11][10] ,
         \registers[11][9] , \registers[11][8] , \registers[11][7] ,
         \registers[11][6] , \registers[11][5] , \registers[11][4] ,
         \registers[11][3] , \registers[11][2] , \registers[11][1] ,
         \registers[11][0] , \registers[12][31] , \registers[12][30] ,
         \registers[12][29] , \registers[12][28] , \registers[12][27] ,
         \registers[12][26] , \registers[12][25] , \registers[12][24] ,
         \registers[12][23] , \registers[12][22] , \registers[12][21] ,
         \registers[12][20] , \registers[12][19] , \registers[12][18] ,
         \registers[12][17] , \registers[12][16] , \registers[12][15] ,
         \registers[12][14] , \registers[12][13] , \registers[12][12] ,
         \registers[12][11] , \registers[12][10] , \registers[12][9] ,
         \registers[12][8] , \registers[12][7] , \registers[12][6] ,
         \registers[12][5] , \registers[12][4] , \registers[12][3] ,
         \registers[12][2] , \registers[12][1] , \registers[12][0] ,
         \registers[13][31] , \registers[13][30] , \registers[13][29] ,
         \registers[13][28] , \registers[13][27] , \registers[13][26] ,
         \registers[13][25] , \registers[13][24] , \registers[13][23] ,
         \registers[13][22] , \registers[13][21] , \registers[13][20] ,
         \registers[13][19] , \registers[13][18] , \registers[13][17] ,
         \registers[13][16] , \registers[13][15] , \registers[13][14] ,
         \registers[13][13] , \registers[13][12] , \registers[13][11] ,
         \registers[13][10] , \registers[13][9] , \registers[13][8] ,
         \registers[13][7] , \registers[13][6] , \registers[13][5] ,
         \registers[13][4] , \registers[13][3] , \registers[13][2] ,
         \registers[13][1] , \registers[13][0] , \registers[14][31] ,
         \registers[14][30] , \registers[14][29] , \registers[14][28] ,
         \registers[14][27] , \registers[14][26] , \registers[14][25] ,
         \registers[14][24] , \registers[14][23] , \registers[14][22] ,
         \registers[14][21] , \registers[14][20] , \registers[14][19] ,
         \registers[14][18] , \registers[14][17] , \registers[14][16] ,
         \registers[14][15] , \registers[14][14] , \registers[14][13] ,
         \registers[14][12] , \registers[14][11] , \registers[14][10] ,
         \registers[14][9] , \registers[14][8] , \registers[14][7] ,
         \registers[14][6] , \registers[14][5] , \registers[14][4] ,
         \registers[14][3] , \registers[14][2] , \registers[14][1] ,
         \registers[14][0] , \registers[15][31] , \registers[15][30] ,
         \registers[15][29] , \registers[15][28] , \registers[15][27] ,
         \registers[15][26] , \registers[15][25] , \registers[15][24] ,
         \registers[15][23] , \registers[15][22] , \registers[15][21] ,
         \registers[15][20] , \registers[15][19] , \registers[15][18] ,
         \registers[15][17] , \registers[15][16] , \registers[15][15] ,
         \registers[15][14] , \registers[15][13] , \registers[15][12] ,
         \registers[15][11] , \registers[15][10] , \registers[15][9] ,
         \registers[15][8] , \registers[15][7] , \registers[15][6] ,
         \registers[15][5] , \registers[15][4] , \registers[15][3] ,
         \registers[15][2] , \registers[15][1] , \registers[15][0] ,
         \registers[16][31] , \registers[16][30] , \registers[16][29] ,
         \registers[16][28] , \registers[16][27] , \registers[16][26] ,
         \registers[16][25] , \registers[16][24] , \registers[16][23] ,
         \registers[16][22] , \registers[16][21] , \registers[16][20] ,
         \registers[16][19] , \registers[16][18] , \registers[16][17] ,
         \registers[16][16] , \registers[16][15] , \registers[16][14] ,
         \registers[16][13] , \registers[16][12] , \registers[16][11] ,
         \registers[16][10] , \registers[16][9] , \registers[16][8] ,
         \registers[16][7] , \registers[16][6] , \registers[16][5] ,
         \registers[16][4] , \registers[16][3] , \registers[16][2] ,
         \registers[16][1] , \registers[16][0] , \registers[17][31] ,
         \registers[17][30] , \registers[17][29] , \registers[17][28] ,
         \registers[17][27] , \registers[17][26] , \registers[17][25] ,
         \registers[17][24] , \registers[17][23] , \registers[17][22] ,
         \registers[17][21] , \registers[17][20] , \registers[17][19] ,
         \registers[17][18] , \registers[17][17] , \registers[17][16] ,
         \registers[17][15] , \registers[17][14] , \registers[17][13] ,
         \registers[17][12] , \registers[17][11] , \registers[17][10] ,
         \registers[17][9] , \registers[17][8] , \registers[17][7] ,
         \registers[17][6] , \registers[17][5] , \registers[17][4] ,
         \registers[17][3] , \registers[17][2] , \registers[17][1] ,
         \registers[17][0] , \registers[18][31] , \registers[18][30] ,
         \registers[18][29] , \registers[18][28] , \registers[18][27] ,
         \registers[18][26] , \registers[18][25] , \registers[18][24] ,
         \registers[18][23] , \registers[18][22] , \registers[18][21] ,
         \registers[18][20] , \registers[18][19] , \registers[18][18] ,
         \registers[18][17] , \registers[18][16] , \registers[18][15] ,
         \registers[18][14] , \registers[18][13] , \registers[18][12] ,
         \registers[18][11] , \registers[18][10] , \registers[18][9] ,
         \registers[18][8] , \registers[18][7] , \registers[18][6] ,
         \registers[18][5] , \registers[18][4] , \registers[18][3] ,
         \registers[18][2] , \registers[18][1] , \registers[18][0] ,
         \registers[19][31] , \registers[19][30] , \registers[19][29] ,
         \registers[19][28] , \registers[19][27] , \registers[19][26] ,
         \registers[19][25] , \registers[19][24] , \registers[19][23] ,
         \registers[19][22] , \registers[19][21] , \registers[19][20] ,
         \registers[19][19] , \registers[19][18] , \registers[19][17] ,
         \registers[19][16] , \registers[19][15] , \registers[19][14] ,
         \registers[19][13] , \registers[19][12] , \registers[19][11] ,
         \registers[19][10] , \registers[19][9] , \registers[19][8] ,
         \registers[19][7] , \registers[19][6] , \registers[19][5] ,
         \registers[19][4] , \registers[19][3] , \registers[19][2] ,
         \registers[19][1] , \registers[19][0] , \registers[20][31] ,
         \registers[20][30] , \registers[20][29] , \registers[20][28] ,
         \registers[20][27] , \registers[20][26] , \registers[20][25] ,
         \registers[20][24] , \registers[20][23] , \registers[20][22] ,
         \registers[20][21] , \registers[20][20] , \registers[20][19] ,
         \registers[20][18] , \registers[20][17] , \registers[20][16] ,
         \registers[20][15] , \registers[20][14] , \registers[20][13] ,
         \registers[20][12] , \registers[20][11] , \registers[20][10] ,
         \registers[20][9] , \registers[20][8] , \registers[20][7] ,
         \registers[20][6] , \registers[20][5] , \registers[20][4] ,
         \registers[20][3] , \registers[20][2] , \registers[20][1] ,
         \registers[20][0] , \registers[21][31] , \registers[21][30] ,
         \registers[21][29] , \registers[21][28] , \registers[21][27] ,
         \registers[21][26] , \registers[21][25] , \registers[21][24] ,
         \registers[21][23] , \registers[21][22] , \registers[21][21] ,
         \registers[21][20] , \registers[21][19] , \registers[21][18] ,
         \registers[21][17] , \registers[21][16] , \registers[21][15] ,
         \registers[21][14] , \registers[21][13] , \registers[21][12] ,
         \registers[21][11] , \registers[21][10] , \registers[21][9] ,
         \registers[21][8] , \registers[21][7] , \registers[21][6] ,
         \registers[21][5] , \registers[21][4] , \registers[21][3] ,
         \registers[21][2] , \registers[21][1] , \registers[21][0] ,
         \registers[22][31] , \registers[22][30] , \registers[22][29] ,
         \registers[22][28] , \registers[22][27] , \registers[22][26] ,
         \registers[22][25] , \registers[22][24] , \registers[22][23] ,
         \registers[22][22] , \registers[22][21] , \registers[22][20] ,
         \registers[22][19] , \registers[22][18] , \registers[22][17] ,
         \registers[22][16] , \registers[22][15] , \registers[22][14] ,
         \registers[22][13] , \registers[22][12] , \registers[22][11] ,
         \registers[22][10] , \registers[22][9] , \registers[22][8] ,
         \registers[22][7] , \registers[22][6] , \registers[22][5] ,
         \registers[22][4] , \registers[22][3] , \registers[22][2] ,
         \registers[22][1] , \registers[22][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[24][31] , \registers[24][30] ,
         \registers[24][29] , \registers[24][28] , \registers[24][27] ,
         \registers[24][26] , \registers[24][25] , \registers[24][24] ,
         \registers[24][23] , \registers[24][22] , \registers[24][21] ,
         \registers[24][20] , \registers[24][19] , \registers[24][18] ,
         \registers[24][17] , \registers[24][16] , \registers[24][15] ,
         \registers[24][14] , \registers[24][13] , \registers[24][12] ,
         \registers[24][11] , \registers[24][10] , \registers[24][9] ,
         \registers[24][8] , \registers[24][7] , \registers[24][6] ,
         \registers[24][5] , \registers[24][4] , \registers[24][3] ,
         \registers[24][2] , \registers[24][1] , \registers[24][0] ,
         \registers[25][31] , \registers[25][30] , \registers[25][29] ,
         \registers[25][28] , \registers[25][27] , \registers[25][26] ,
         \registers[25][25] , \registers[25][24] , \registers[25][23] ,
         \registers[25][22] , \registers[25][21] , \registers[25][20] ,
         \registers[25][19] , \registers[25][18] , \registers[25][17] ,
         \registers[25][16] , \registers[25][15] , \registers[25][14] ,
         \registers[25][13] , \registers[25][12] , \registers[25][11] ,
         \registers[25][10] , \registers[25][9] , \registers[25][8] ,
         \registers[25][7] , \registers[25][6] , \registers[25][5] ,
         \registers[25][4] , \registers[25][3] , \registers[25][2] ,
         \registers[25][1] , \registers[25][0] , \registers[26][31] ,
         \registers[26][30] , \registers[26][29] , \registers[26][28] ,
         \registers[26][27] , \registers[26][26] , \registers[26][25] ,
         \registers[26][24] , \registers[26][23] , \registers[26][22] ,
         \registers[26][21] , \registers[26][20] , \registers[26][19] ,
         \registers[26][18] , \registers[26][17] , \registers[26][16] ,
         \registers[26][15] , \registers[26][14] , \registers[26][13] ,
         \registers[26][12] , \registers[26][11] , \registers[26][10] ,
         \registers[26][9] , \registers[26][8] , \registers[26][7] ,
         \registers[26][6] , \registers[26][5] , \registers[26][4] ,
         \registers[26][3] , \registers[26][2] , \registers[26][1] ,
         \registers[26][0] , \registers[27][31] , \registers[27][30] ,
         \registers[27][29] , \registers[27][28] , \registers[27][27] ,
         \registers[27][26] , \registers[27][25] , \registers[27][24] ,
         \registers[27][23] , \registers[27][22] , \registers[27][21] ,
         \registers[27][20] , \registers[27][19] , \registers[27][18] ,
         \registers[27][17] , \registers[27][16] , \registers[27][15] ,
         \registers[27][14] , \registers[27][13] , \registers[27][12] ,
         \registers[27][11] , \registers[27][10] , \registers[27][9] ,
         \registers[27][8] , \registers[27][7] , \registers[27][6] ,
         \registers[27][5] , \registers[27][4] , \registers[27][3] ,
         \registers[27][2] , \registers[27][1] , \registers[27][0] ,
         \registers[28][31] , \registers[28][30] , \registers[28][29] ,
         \registers[28][28] , \registers[28][27] , \registers[28][26] ,
         \registers[28][25] , \registers[28][24] , \registers[28][23] ,
         \registers[28][22] , \registers[28][21] , \registers[28][20] ,
         \registers[28][19] , \registers[28][18] , \registers[28][17] ,
         \registers[28][16] , \registers[28][15] , \registers[28][14] ,
         \registers[28][13] , \registers[28][12] , \registers[28][11] ,
         \registers[28][10] , \registers[28][9] , \registers[28][8] ,
         \registers[28][7] , \registers[28][6] , \registers[28][5] ,
         \registers[28][4] , \registers[28][3] , \registers[28][2] ,
         \registers[28][1] , \registers[28][0] , \registers[29][31] ,
         \registers[29][30] , \registers[29][29] , \registers[29][28] ,
         \registers[29][27] , \registers[29][26] , \registers[29][25] ,
         \registers[29][24] , \registers[29][23] , \registers[29][22] ,
         \registers[29][21] , \registers[29][20] , \registers[29][19] ,
         \registers[29][18] , \registers[29][17] , \registers[29][16] ,
         \registers[29][15] , \registers[29][14] , \registers[29][13] ,
         \registers[29][12] , \registers[29][11] , \registers[29][10] ,
         \registers[29][9] , \registers[29][8] , \registers[29][7] ,
         \registers[29][6] , \registers[29][5] , \registers[29][4] ,
         \registers[29][3] , \registers[29][2] , \registers[29][1] ,
         \registers[29][0] , \registers[30][31] , \registers[30][30] ,
         \registers[30][29] , \registers[30][28] , \registers[30][27] ,
         \registers[30][26] , \registers[30][25] , \registers[30][24] ,
         \registers[30][23] , \registers[30][22] , \registers[30][21] ,
         \registers[30][20] , \registers[30][19] , \registers[30][18] ,
         \registers[30][17] , \registers[30][16] , \registers[30][15] ,
         \registers[30][14] , \registers[30][13] , \registers[30][12] ,
         \registers[30][11] , \registers[30][10] , \registers[30][9] ,
         \registers[30][8] , \registers[30][7] , \registers[30][6] ,
         \registers[30][5] , \registers[30][4] , \registers[30][3] ,
         \registers[30][2] , \registers[30][1] , \registers[30][0] ,
         \registers[31][31] , \registers[31][30] , \registers[31][29] ,
         \registers[31][28] , \registers[31][27] , \registers[31][26] ,
         \registers[31][25] , \registers[31][24] , \registers[31][23] ,
         \registers[31][22] , \registers[31][21] , \registers[31][20] ,
         \registers[31][19] , \registers[31][18] , \registers[31][17] ,
         \registers[31][16] , \registers[31][15] , \registers[31][14] ,
         \registers[31][13] , \registers[31][12] , \registers[31][11] ,
         \registers[31][10] , \registers[31][9] , \registers[31][8] ,
         \registers[31][7] , \registers[31][6] , \registers[31][5] ,
         \registers[31][4] , \registers[31][3] , \registers[31][2] ,
         \registers[31][1] , \registers[31][0] , N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N243, N244, N245, N246, N247, N248,
         N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N307, N308, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
         N369, N371, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689;

  DLH_X1 \registers_reg[1][31]  ( .G(n1970), .D(n2060), .Q(\registers[1][31] )
         );
  DLH_X1 \registers_reg[1][30]  ( .G(n1970), .D(n2063), .Q(\registers[1][30] )
         );
  DLH_X1 \registers_reg[1][29]  ( .G(n1970), .D(n2066), .Q(\registers[1][29] )
         );
  DLH_X1 \registers_reg[1][28]  ( .G(n1970), .D(n2069), .Q(\registers[1][28] )
         );
  DLH_X1 \registers_reg[1][27]  ( .G(n1970), .D(n2072), .Q(\registers[1][27] )
         );
  DLH_X1 \registers_reg[1][26]  ( .G(n1970), .D(n2075), .Q(\registers[1][26] )
         );
  DLH_X1 \registers_reg[1][25]  ( .G(n1970), .D(n2078), .Q(\registers[1][25] )
         );
  DLH_X1 \registers_reg[1][24]  ( .G(n1969), .D(n2081), .Q(\registers[1][24] )
         );
  DLH_X1 \registers_reg[1][23]  ( .G(n1969), .D(n2084), .Q(\registers[1][23] )
         );
  DLH_X1 \registers_reg[1][22]  ( .G(n1969), .D(n2087), .Q(\registers[1][22] )
         );
  DLH_X1 \registers_reg[1][21]  ( .G(n1969), .D(n2090), .Q(\registers[1][21] )
         );
  DLH_X1 \registers_reg[1][20]  ( .G(n1970), .D(n2093), .Q(\registers[1][20] )
         );
  DLH_X1 \registers_reg[1][19]  ( .G(n1969), .D(n2096), .Q(\registers[1][19] )
         );
  DLH_X1 \registers_reg[1][18]  ( .G(n1969), .D(n2099), .Q(\registers[1][18] )
         );
  DLH_X1 \registers_reg[1][17]  ( .G(n1970), .D(n2102), .Q(\registers[1][17] )
         );
  DLH_X1 \registers_reg[1][16]  ( .G(n1969), .D(n2105), .Q(\registers[1][16] )
         );
  DLH_X1 \registers_reg[1][15]  ( .G(n1969), .D(n2108), .Q(\registers[1][15] )
         );
  DLH_X1 \registers_reg[1][14]  ( .G(n1969), .D(n2111), .Q(\registers[1][14] )
         );
  DLH_X1 \registers_reg[1][13]  ( .G(n1968), .D(n2114), .Q(\registers[1][13] )
         );
  DLH_X1 \registers_reg[1][12]  ( .G(n1969), .D(n2117), .Q(\registers[1][12] )
         );
  DLH_X1 \registers_reg[1][11]  ( .G(n1968), .D(n2120), .Q(\registers[1][11] )
         );
  DLH_X1 \registers_reg[1][10]  ( .G(n1968), .D(n2123), .Q(\registers[1][10] )
         );
  DLH_X1 \registers_reg[1][9]  ( .G(n1968), .D(n2126), .Q(\registers[1][9] )
         );
  DLH_X1 \registers_reg[1][8]  ( .G(n1968), .D(n2129), .Q(\registers[1][8] )
         );
  DLH_X1 \registers_reg[1][7]  ( .G(n1968), .D(n2132), .Q(\registers[1][7] )
         );
  DLH_X1 \registers_reg[1][6]  ( .G(n1968), .D(n2135), .Q(\registers[1][6] )
         );
  DLH_X1 \registers_reg[1][5]  ( .G(n1968), .D(n2138), .Q(\registers[1][5] )
         );
  DLH_X1 \registers_reg[1][4]  ( .G(n1968), .D(n2141), .Q(\registers[1][4] )
         );
  DLH_X1 \registers_reg[1][3]  ( .G(n1968), .D(n2144), .Q(\registers[1][3] )
         );
  DLH_X1 \registers_reg[1][2]  ( .G(n1968), .D(n2147), .Q(\registers[1][2] )
         );
  DLH_X1 \registers_reg[1][1]  ( .G(n1969), .D(n2150), .Q(\registers[1][1] )
         );
  DLH_X1 \registers_reg[1][0]  ( .G(n1970), .D(n2153), .Q(\registers[1][0] )
         );
  DLH_X1 \registers_reg[2][31]  ( .G(n1973), .D(n2060), .Q(\registers[2][31] )
         );
  DLH_X1 \registers_reg[2][30]  ( .G(n1973), .D(n2063), .Q(\registers[2][30] )
         );
  DLH_X1 \registers_reg[2][29]  ( .G(n1973), .D(n2066), .Q(\registers[2][29] )
         );
  DLH_X1 \registers_reg[2][28]  ( .G(n1973), .D(n2069), .Q(\registers[2][28] )
         );
  DLH_X1 \registers_reg[2][27]  ( .G(n1973), .D(n2072), .Q(\registers[2][27] )
         );
  DLH_X1 \registers_reg[2][26]  ( .G(n1973), .D(n2075), .Q(\registers[2][26] )
         );
  DLH_X1 \registers_reg[2][25]  ( .G(n1973), .D(n2078), .Q(\registers[2][25] )
         );
  DLH_X1 \registers_reg[2][24]  ( .G(n1972), .D(n2081), .Q(\registers[2][24] )
         );
  DLH_X1 \registers_reg[2][23]  ( .G(n1972), .D(n2084), .Q(\registers[2][23] )
         );
  DLH_X1 \registers_reg[2][22]  ( .G(n1972), .D(n2087), .Q(\registers[2][22] )
         );
  DLH_X1 \registers_reg[2][21]  ( .G(n1972), .D(n2090), .Q(\registers[2][21] )
         );
  DLH_X1 \registers_reg[2][20]  ( .G(n1973), .D(n2093), .Q(\registers[2][20] )
         );
  DLH_X1 \registers_reg[2][19]  ( .G(n1972), .D(n2096), .Q(\registers[2][19] )
         );
  DLH_X1 \registers_reg[2][18]  ( .G(n1972), .D(n2099), .Q(\registers[2][18] )
         );
  DLH_X1 \registers_reg[2][17]  ( .G(n1973), .D(n2102), .Q(\registers[2][17] )
         );
  DLH_X1 \registers_reg[2][16]  ( .G(n1972), .D(n2105), .Q(\registers[2][16] )
         );
  DLH_X1 \registers_reg[2][15]  ( .G(n1972), .D(n2108), .Q(\registers[2][15] )
         );
  DLH_X1 \registers_reg[2][14]  ( .G(n1972), .D(n2111), .Q(\registers[2][14] )
         );
  DLH_X1 \registers_reg[2][13]  ( .G(n1971), .D(n2114), .Q(\registers[2][13] )
         );
  DLH_X1 \registers_reg[2][12]  ( .G(n1972), .D(n2117), .Q(\registers[2][12] )
         );
  DLH_X1 \registers_reg[2][11]  ( .G(n1971), .D(n2120), .Q(\registers[2][11] )
         );
  DLH_X1 \registers_reg[2][10]  ( .G(n1971), .D(n2123), .Q(\registers[2][10] )
         );
  DLH_X1 \registers_reg[2][9]  ( .G(n1971), .D(n2126), .Q(\registers[2][9] )
         );
  DLH_X1 \registers_reg[2][8]  ( .G(n1971), .D(n2129), .Q(\registers[2][8] )
         );
  DLH_X1 \registers_reg[2][7]  ( .G(n1971), .D(n2132), .Q(\registers[2][7] )
         );
  DLH_X1 \registers_reg[2][6]  ( .G(n1971), .D(n2135), .Q(\registers[2][6] )
         );
  DLH_X1 \registers_reg[2][5]  ( .G(n1971), .D(n2138), .Q(\registers[2][5] )
         );
  DLH_X1 \registers_reg[2][4]  ( .G(n1971), .D(n2141), .Q(\registers[2][4] )
         );
  DLH_X1 \registers_reg[2][3]  ( .G(n1971), .D(n2144), .Q(\registers[2][3] )
         );
  DLH_X1 \registers_reg[2][2]  ( .G(n1971), .D(n2147), .Q(\registers[2][2] )
         );
  DLH_X1 \registers_reg[2][1]  ( .G(n1972), .D(n2150), .Q(\registers[2][1] )
         );
  DLH_X1 \registers_reg[2][0]  ( .G(n1973), .D(n2153), .Q(\registers[2][0] )
         );
  DLH_X1 \registers_reg[3][31]  ( .G(n1976), .D(n2060), .Q(\registers[3][31] )
         );
  DLH_X1 \registers_reg[3][30]  ( .G(n1976), .D(n2063), .Q(\registers[3][30] )
         );
  DLH_X1 \registers_reg[3][29]  ( .G(n1976), .D(n2066), .Q(\registers[3][29] )
         );
  DLH_X1 \registers_reg[3][28]  ( .G(n1976), .D(n2069), .Q(\registers[3][28] )
         );
  DLH_X1 \registers_reg[3][27]  ( .G(n1976), .D(n2072), .Q(\registers[3][27] )
         );
  DLH_X1 \registers_reg[3][26]  ( .G(n1976), .D(n2075), .Q(\registers[3][26] )
         );
  DLH_X1 \registers_reg[3][25]  ( .G(n1976), .D(n2078), .Q(\registers[3][25] )
         );
  DLH_X1 \registers_reg[3][24]  ( .G(n1975), .D(n2081), .Q(\registers[3][24] )
         );
  DLH_X1 \registers_reg[3][23]  ( .G(n1975), .D(n2084), .Q(\registers[3][23] )
         );
  DLH_X1 \registers_reg[3][22]  ( .G(n1975), .D(n2087), .Q(\registers[3][22] )
         );
  DLH_X1 \registers_reg[3][21]  ( .G(n1975), .D(n2090), .Q(\registers[3][21] )
         );
  DLH_X1 \registers_reg[3][20]  ( .G(n1976), .D(n2093), .Q(\registers[3][20] )
         );
  DLH_X1 \registers_reg[3][19]  ( .G(n1975), .D(n2096), .Q(\registers[3][19] )
         );
  DLH_X1 \registers_reg[3][18]  ( .G(n1975), .D(n2099), .Q(\registers[3][18] )
         );
  DLH_X1 \registers_reg[3][17]  ( .G(n1976), .D(n2102), .Q(\registers[3][17] )
         );
  DLH_X1 \registers_reg[3][16]  ( .G(n1975), .D(n2105), .Q(\registers[3][16] )
         );
  DLH_X1 \registers_reg[3][15]  ( .G(n1975), .D(n2108), .Q(\registers[3][15] )
         );
  DLH_X1 \registers_reg[3][14]  ( .G(n1975), .D(n2111), .Q(\registers[3][14] )
         );
  DLH_X1 \registers_reg[3][13]  ( .G(n1974), .D(n2114), .Q(\registers[3][13] )
         );
  DLH_X1 \registers_reg[3][12]  ( .G(n1975), .D(n2117), .Q(\registers[3][12] )
         );
  DLH_X1 \registers_reg[3][11]  ( .G(n1974), .D(n2120), .Q(\registers[3][11] )
         );
  DLH_X1 \registers_reg[3][10]  ( .G(n1974), .D(n2123), .Q(\registers[3][10] )
         );
  DLH_X1 \registers_reg[3][9]  ( .G(n1974), .D(n2126), .Q(\registers[3][9] )
         );
  DLH_X1 \registers_reg[3][8]  ( .G(n1974), .D(n2129), .Q(\registers[3][8] )
         );
  DLH_X1 \registers_reg[3][7]  ( .G(n1974), .D(n2132), .Q(\registers[3][7] )
         );
  DLH_X1 \registers_reg[3][6]  ( .G(n1974), .D(n2135), .Q(\registers[3][6] )
         );
  DLH_X1 \registers_reg[3][5]  ( .G(n1974), .D(n2138), .Q(\registers[3][5] )
         );
  DLH_X1 \registers_reg[3][4]  ( .G(n1974), .D(n2141), .Q(\registers[3][4] )
         );
  DLH_X1 \registers_reg[3][3]  ( .G(n1974), .D(n2144), .Q(\registers[3][3] )
         );
  DLH_X1 \registers_reg[3][2]  ( .G(n1974), .D(n2147), .Q(\registers[3][2] )
         );
  DLH_X1 \registers_reg[3][1]  ( .G(n1975), .D(n2150), .Q(\registers[3][1] )
         );
  DLH_X1 \registers_reg[3][0]  ( .G(n1976), .D(n2153), .Q(\registers[3][0] )
         );
  DLH_X1 \registers_reg[4][31]  ( .G(n1979), .D(n2060), .Q(\registers[4][31] )
         );
  DLH_X1 \registers_reg[4][30]  ( .G(n1979), .D(n2063), .Q(\registers[4][30] )
         );
  DLH_X1 \registers_reg[4][29]  ( .G(n1979), .D(n2066), .Q(\registers[4][29] )
         );
  DLH_X1 \registers_reg[4][28]  ( .G(n1979), .D(n2069), .Q(\registers[4][28] )
         );
  DLH_X1 \registers_reg[4][27]  ( .G(n1979), .D(n2072), .Q(\registers[4][27] )
         );
  DLH_X1 \registers_reg[4][26]  ( .G(n1979), .D(n2075), .Q(\registers[4][26] )
         );
  DLH_X1 \registers_reg[4][25]  ( .G(n1979), .D(n2078), .Q(\registers[4][25] )
         );
  DLH_X1 \registers_reg[4][24]  ( .G(n1978), .D(n2081), .Q(\registers[4][24] )
         );
  DLH_X1 \registers_reg[4][23]  ( .G(n1978), .D(n2084), .Q(\registers[4][23] )
         );
  DLH_X1 \registers_reg[4][22]  ( .G(n1978), .D(n2087), .Q(\registers[4][22] )
         );
  DLH_X1 \registers_reg[4][21]  ( .G(n1978), .D(n2090), .Q(\registers[4][21] )
         );
  DLH_X1 \registers_reg[4][20]  ( .G(n1979), .D(n2093), .Q(\registers[4][20] )
         );
  DLH_X1 \registers_reg[4][19]  ( .G(n1978), .D(n2096), .Q(\registers[4][19] )
         );
  DLH_X1 \registers_reg[4][18]  ( .G(n1978), .D(n2099), .Q(\registers[4][18] )
         );
  DLH_X1 \registers_reg[4][17]  ( .G(n1979), .D(n2102), .Q(\registers[4][17] )
         );
  DLH_X1 \registers_reg[4][16]  ( .G(n1978), .D(n2105), .Q(\registers[4][16] )
         );
  DLH_X1 \registers_reg[4][15]  ( .G(n1978), .D(n2108), .Q(\registers[4][15] )
         );
  DLH_X1 \registers_reg[4][14]  ( .G(n1978), .D(n2111), .Q(\registers[4][14] )
         );
  DLH_X1 \registers_reg[4][13]  ( .G(n1977), .D(n2114), .Q(\registers[4][13] )
         );
  DLH_X1 \registers_reg[4][12]  ( .G(n1978), .D(n2117), .Q(\registers[4][12] )
         );
  DLH_X1 \registers_reg[4][11]  ( .G(n1977), .D(n2120), .Q(\registers[4][11] )
         );
  DLH_X1 \registers_reg[4][10]  ( .G(n1977), .D(n2123), .Q(\registers[4][10] )
         );
  DLH_X1 \registers_reg[4][9]  ( .G(n1977), .D(n2126), .Q(\registers[4][9] )
         );
  DLH_X1 \registers_reg[4][8]  ( .G(n1977), .D(n2129), .Q(\registers[4][8] )
         );
  DLH_X1 \registers_reg[4][7]  ( .G(n1977), .D(n2132), .Q(\registers[4][7] )
         );
  DLH_X1 \registers_reg[4][6]  ( .G(n1977), .D(n2135), .Q(\registers[4][6] )
         );
  DLH_X1 \registers_reg[4][5]  ( .G(n1977), .D(n2138), .Q(\registers[4][5] )
         );
  DLH_X1 \registers_reg[4][4]  ( .G(n1977), .D(n2141), .Q(\registers[4][4] )
         );
  DLH_X1 \registers_reg[4][3]  ( .G(n1977), .D(n2144), .Q(\registers[4][3] )
         );
  DLH_X1 \registers_reg[4][2]  ( .G(n1977), .D(n2147), .Q(\registers[4][2] )
         );
  DLH_X1 \registers_reg[4][1]  ( .G(n1978), .D(n2150), .Q(\registers[4][1] )
         );
  DLH_X1 \registers_reg[4][0]  ( .G(n1979), .D(n2153), .Q(\registers[4][0] )
         );
  DLH_X1 \registers_reg[5][31]  ( .G(n1982), .D(n2060), .Q(\registers[5][31] )
         );
  DLH_X1 \registers_reg[5][30]  ( .G(n1982), .D(n2063), .Q(\registers[5][30] )
         );
  DLH_X1 \registers_reg[5][29]  ( .G(n1982), .D(n2066), .Q(\registers[5][29] )
         );
  DLH_X1 \registers_reg[5][28]  ( .G(n1982), .D(n2069), .Q(\registers[5][28] )
         );
  DLH_X1 \registers_reg[5][27]  ( .G(n1982), .D(n2072), .Q(\registers[5][27] )
         );
  DLH_X1 \registers_reg[5][26]  ( .G(n1982), .D(n2075), .Q(\registers[5][26] )
         );
  DLH_X1 \registers_reg[5][25]  ( .G(n1982), .D(n2078), .Q(\registers[5][25] )
         );
  DLH_X1 \registers_reg[5][24]  ( .G(n1981), .D(n2081), .Q(\registers[5][24] )
         );
  DLH_X1 \registers_reg[5][23]  ( .G(n1981), .D(n2084), .Q(\registers[5][23] )
         );
  DLH_X1 \registers_reg[5][22]  ( .G(n1981), .D(n2087), .Q(\registers[5][22] )
         );
  DLH_X1 \registers_reg[5][21]  ( .G(n1981), .D(n2090), .Q(\registers[5][21] )
         );
  DLH_X1 \registers_reg[5][20]  ( .G(n1982), .D(n2093), .Q(\registers[5][20] )
         );
  DLH_X1 \registers_reg[5][19]  ( .G(n1981), .D(n2096), .Q(\registers[5][19] )
         );
  DLH_X1 \registers_reg[5][18]  ( .G(n1981), .D(n2099), .Q(\registers[5][18] )
         );
  DLH_X1 \registers_reg[5][17]  ( .G(n1982), .D(n2102), .Q(\registers[5][17] )
         );
  DLH_X1 \registers_reg[5][16]  ( .G(n1981), .D(n2105), .Q(\registers[5][16] )
         );
  DLH_X1 \registers_reg[5][15]  ( .G(n1981), .D(n2108), .Q(\registers[5][15] )
         );
  DLH_X1 \registers_reg[5][14]  ( .G(n1981), .D(n2111), .Q(\registers[5][14] )
         );
  DLH_X1 \registers_reg[5][13]  ( .G(n1980), .D(n2114), .Q(\registers[5][13] )
         );
  DLH_X1 \registers_reg[5][12]  ( .G(n1981), .D(n2117), .Q(\registers[5][12] )
         );
  DLH_X1 \registers_reg[5][11]  ( .G(n1980), .D(n2120), .Q(\registers[5][11] )
         );
  DLH_X1 \registers_reg[5][10]  ( .G(n1980), .D(n2123), .Q(\registers[5][10] )
         );
  DLH_X1 \registers_reg[5][9]  ( .G(n1980), .D(n2126), .Q(\registers[5][9] )
         );
  DLH_X1 \registers_reg[5][8]  ( .G(n1980), .D(n2129), .Q(\registers[5][8] )
         );
  DLH_X1 \registers_reg[5][7]  ( .G(n1980), .D(n2132), .Q(\registers[5][7] )
         );
  DLH_X1 \registers_reg[5][6]  ( .G(n1980), .D(n2135), .Q(\registers[5][6] )
         );
  DLH_X1 \registers_reg[5][5]  ( .G(n1980), .D(n2138), .Q(\registers[5][5] )
         );
  DLH_X1 \registers_reg[5][4]  ( .G(n1980), .D(n2141), .Q(\registers[5][4] )
         );
  DLH_X1 \registers_reg[5][3]  ( .G(n1980), .D(n2144), .Q(\registers[5][3] )
         );
  DLH_X1 \registers_reg[5][2]  ( .G(n1980), .D(n2147), .Q(\registers[5][2] )
         );
  DLH_X1 \registers_reg[5][1]  ( .G(n1981), .D(n2150), .Q(\registers[5][1] )
         );
  DLH_X1 \registers_reg[5][0]  ( .G(n1982), .D(n2153), .Q(\registers[5][0] )
         );
  DLH_X1 \registers_reg[6][31]  ( .G(n1985), .D(n2060), .Q(\registers[6][31] )
         );
  DLH_X1 \registers_reg[6][30]  ( .G(n1985), .D(n2063), .Q(\registers[6][30] )
         );
  DLH_X1 \registers_reg[6][29]  ( .G(n1985), .D(n2066), .Q(\registers[6][29] )
         );
  DLH_X1 \registers_reg[6][28]  ( .G(n1985), .D(n2069), .Q(\registers[6][28] )
         );
  DLH_X1 \registers_reg[6][27]  ( .G(n1985), .D(n2072), .Q(\registers[6][27] )
         );
  DLH_X1 \registers_reg[6][26]  ( .G(n1985), .D(n2075), .Q(\registers[6][26] )
         );
  DLH_X1 \registers_reg[6][25]  ( .G(n1985), .D(n2078), .Q(\registers[6][25] )
         );
  DLH_X1 \registers_reg[6][24]  ( .G(n1984), .D(n2081), .Q(\registers[6][24] )
         );
  DLH_X1 \registers_reg[6][23]  ( .G(n1984), .D(n2084), .Q(\registers[6][23] )
         );
  DLH_X1 \registers_reg[6][22]  ( .G(n1984), .D(n2087), .Q(\registers[6][22] )
         );
  DLH_X1 \registers_reg[6][21]  ( .G(n1984), .D(n2090), .Q(\registers[6][21] )
         );
  DLH_X1 \registers_reg[6][20]  ( .G(n1985), .D(n2093), .Q(\registers[6][20] )
         );
  DLH_X1 \registers_reg[6][19]  ( .G(n1984), .D(n2096), .Q(\registers[6][19] )
         );
  DLH_X1 \registers_reg[6][18]  ( .G(n1984), .D(n2099), .Q(\registers[6][18] )
         );
  DLH_X1 \registers_reg[6][17]  ( .G(n1985), .D(n2102), .Q(\registers[6][17] )
         );
  DLH_X1 \registers_reg[6][16]  ( .G(n1984), .D(n2105), .Q(\registers[6][16] )
         );
  DLH_X1 \registers_reg[6][15]  ( .G(n1984), .D(n2108), .Q(\registers[6][15] )
         );
  DLH_X1 \registers_reg[6][14]  ( .G(n1984), .D(n2111), .Q(\registers[6][14] )
         );
  DLH_X1 \registers_reg[6][13]  ( .G(n1983), .D(n2114), .Q(\registers[6][13] )
         );
  DLH_X1 \registers_reg[6][12]  ( .G(n1984), .D(n2117), .Q(\registers[6][12] )
         );
  DLH_X1 \registers_reg[6][11]  ( .G(n1983), .D(n2120), .Q(\registers[6][11] )
         );
  DLH_X1 \registers_reg[6][10]  ( .G(n1983), .D(n2123), .Q(\registers[6][10] )
         );
  DLH_X1 \registers_reg[6][9]  ( .G(n1983), .D(n2126), .Q(\registers[6][9] )
         );
  DLH_X1 \registers_reg[6][8]  ( .G(n1983), .D(n2129), .Q(\registers[6][8] )
         );
  DLH_X1 \registers_reg[6][7]  ( .G(n1983), .D(n2132), .Q(\registers[6][7] )
         );
  DLH_X1 \registers_reg[6][6]  ( .G(n1983), .D(n2135), .Q(\registers[6][6] )
         );
  DLH_X1 \registers_reg[6][5]  ( .G(n1983), .D(n2138), .Q(\registers[6][5] )
         );
  DLH_X1 \registers_reg[6][4]  ( .G(n1983), .D(n2141), .Q(\registers[6][4] )
         );
  DLH_X1 \registers_reg[6][3]  ( .G(n1983), .D(n2144), .Q(\registers[6][3] )
         );
  DLH_X1 \registers_reg[6][2]  ( .G(n1983), .D(n2147), .Q(\registers[6][2] )
         );
  DLH_X1 \registers_reg[6][1]  ( .G(n1984), .D(n2150), .Q(\registers[6][1] )
         );
  DLH_X1 \registers_reg[6][0]  ( .G(n1985), .D(n2153), .Q(\registers[6][0] )
         );
  DLH_X1 \registers_reg[7][31]  ( .G(n1988), .D(n2060), .Q(\registers[7][31] )
         );
  DLH_X1 \registers_reg[7][30]  ( .G(n1988), .D(n2063), .Q(\registers[7][30] )
         );
  DLH_X1 \registers_reg[7][29]  ( .G(n1988), .D(n2066), .Q(\registers[7][29] )
         );
  DLH_X1 \registers_reg[7][28]  ( .G(n1988), .D(n2069), .Q(\registers[7][28] )
         );
  DLH_X1 \registers_reg[7][27]  ( .G(n1988), .D(n2072), .Q(\registers[7][27] )
         );
  DLH_X1 \registers_reg[7][26]  ( .G(n1988), .D(n2075), .Q(\registers[7][26] )
         );
  DLH_X1 \registers_reg[7][25]  ( .G(n1988), .D(n2078), .Q(\registers[7][25] )
         );
  DLH_X1 \registers_reg[7][24]  ( .G(n1987), .D(n2081), .Q(\registers[7][24] )
         );
  DLH_X1 \registers_reg[7][23]  ( .G(n1987), .D(n2084), .Q(\registers[7][23] )
         );
  DLH_X1 \registers_reg[7][22]  ( .G(n1987), .D(n2087), .Q(\registers[7][22] )
         );
  DLH_X1 \registers_reg[7][21]  ( .G(n1987), .D(n2090), .Q(\registers[7][21] )
         );
  DLH_X1 \registers_reg[7][20]  ( .G(n1988), .D(n2093), .Q(\registers[7][20] )
         );
  DLH_X1 \registers_reg[7][19]  ( .G(n1987), .D(n2096), .Q(\registers[7][19] )
         );
  DLH_X1 \registers_reg[7][18]  ( .G(n1987), .D(n2099), .Q(\registers[7][18] )
         );
  DLH_X1 \registers_reg[7][17]  ( .G(n1988), .D(n2102), .Q(\registers[7][17] )
         );
  DLH_X1 \registers_reg[7][16]  ( .G(n1987), .D(n2105), .Q(\registers[7][16] )
         );
  DLH_X1 \registers_reg[7][15]  ( .G(n1987), .D(n2108), .Q(\registers[7][15] )
         );
  DLH_X1 \registers_reg[7][14]  ( .G(n1987), .D(n2111), .Q(\registers[7][14] )
         );
  DLH_X1 \registers_reg[7][13]  ( .G(n1986), .D(n2114), .Q(\registers[7][13] )
         );
  DLH_X1 \registers_reg[7][12]  ( .G(n1987), .D(n2117), .Q(\registers[7][12] )
         );
  DLH_X1 \registers_reg[7][11]  ( .G(n1986), .D(n2120), .Q(\registers[7][11] )
         );
  DLH_X1 \registers_reg[7][10]  ( .G(n1986), .D(n2123), .Q(\registers[7][10] )
         );
  DLH_X1 \registers_reg[7][9]  ( .G(n1986), .D(n2126), .Q(\registers[7][9] )
         );
  DLH_X1 \registers_reg[7][8]  ( .G(n1986), .D(n2129), .Q(\registers[7][8] )
         );
  DLH_X1 \registers_reg[7][7]  ( .G(n1986), .D(n2132), .Q(\registers[7][7] )
         );
  DLH_X1 \registers_reg[7][6]  ( .G(n1986), .D(n2135), .Q(\registers[7][6] )
         );
  DLH_X1 \registers_reg[7][5]  ( .G(n1986), .D(n2138), .Q(\registers[7][5] )
         );
  DLH_X1 \registers_reg[7][4]  ( .G(n1986), .D(n2141), .Q(\registers[7][4] )
         );
  DLH_X1 \registers_reg[7][3]  ( .G(n1986), .D(n2144), .Q(\registers[7][3] )
         );
  DLH_X1 \registers_reg[7][2]  ( .G(n1986), .D(n2147), .Q(\registers[7][2] )
         );
  DLH_X1 \registers_reg[7][1]  ( .G(n1987), .D(n2150), .Q(\registers[7][1] )
         );
  DLH_X1 \registers_reg[7][0]  ( .G(n1988), .D(n2153), .Q(\registers[7][0] )
         );
  DLH_X1 \registers_reg[8][31]  ( .G(n1991), .D(n2060), .Q(\registers[8][31] )
         );
  DLH_X1 \registers_reg[8][30]  ( .G(n1991), .D(n2063), .Q(\registers[8][30] )
         );
  DLH_X1 \registers_reg[8][29]  ( .G(n1991), .D(n2066), .Q(\registers[8][29] )
         );
  DLH_X1 \registers_reg[8][28]  ( .G(n1991), .D(n2069), .Q(\registers[8][28] )
         );
  DLH_X1 \registers_reg[8][27]  ( .G(n1991), .D(n2072), .Q(\registers[8][27] )
         );
  DLH_X1 \registers_reg[8][26]  ( .G(n1991), .D(n2075), .Q(\registers[8][26] )
         );
  DLH_X1 \registers_reg[8][25]  ( .G(n1991), .D(n2078), .Q(\registers[8][25] )
         );
  DLH_X1 \registers_reg[8][24]  ( .G(n1990), .D(n2081), .Q(\registers[8][24] )
         );
  DLH_X1 \registers_reg[8][23]  ( .G(n1990), .D(n2084), .Q(\registers[8][23] )
         );
  DLH_X1 \registers_reg[8][22]  ( .G(n1990), .D(n2087), .Q(\registers[8][22] )
         );
  DLH_X1 \registers_reg[8][21]  ( .G(n1990), .D(n2090), .Q(\registers[8][21] )
         );
  DLH_X1 \registers_reg[8][20]  ( .G(n1991), .D(n2093), .Q(\registers[8][20] )
         );
  DLH_X1 \registers_reg[8][19]  ( .G(n1990), .D(n2096), .Q(\registers[8][19] )
         );
  DLH_X1 \registers_reg[8][18]  ( .G(n1990), .D(n2099), .Q(\registers[8][18] )
         );
  DLH_X1 \registers_reg[8][17]  ( .G(n1991), .D(n2102), .Q(\registers[8][17] )
         );
  DLH_X1 \registers_reg[8][16]  ( .G(n1990), .D(n2105), .Q(\registers[8][16] )
         );
  DLH_X1 \registers_reg[8][15]  ( .G(n1990), .D(n2108), .Q(\registers[8][15] )
         );
  DLH_X1 \registers_reg[8][14]  ( .G(n1990), .D(n2111), .Q(\registers[8][14] )
         );
  DLH_X1 \registers_reg[8][13]  ( .G(n1989), .D(n2114), .Q(\registers[8][13] )
         );
  DLH_X1 \registers_reg[8][12]  ( .G(n1990), .D(n2117), .Q(\registers[8][12] )
         );
  DLH_X1 \registers_reg[8][11]  ( .G(n1989), .D(n2120), .Q(\registers[8][11] )
         );
  DLH_X1 \registers_reg[8][10]  ( .G(n1989), .D(n2123), .Q(\registers[8][10] )
         );
  DLH_X1 \registers_reg[8][9]  ( .G(n1989), .D(n2126), .Q(\registers[8][9] )
         );
  DLH_X1 \registers_reg[8][8]  ( .G(n1989), .D(n2129), .Q(\registers[8][8] )
         );
  DLH_X1 \registers_reg[8][7]  ( .G(n1989), .D(n2132), .Q(\registers[8][7] )
         );
  DLH_X1 \registers_reg[8][6]  ( .G(n1989), .D(n2135), .Q(\registers[8][6] )
         );
  DLH_X1 \registers_reg[8][5]  ( .G(n1989), .D(n2138), .Q(\registers[8][5] )
         );
  DLH_X1 \registers_reg[8][4]  ( .G(n1989), .D(n2141), .Q(\registers[8][4] )
         );
  DLH_X1 \registers_reg[8][3]  ( .G(n1989), .D(n2144), .Q(\registers[8][3] )
         );
  DLH_X1 \registers_reg[8][2]  ( .G(n1989), .D(n2147), .Q(\registers[8][2] )
         );
  DLH_X1 \registers_reg[8][1]  ( .G(n1990), .D(n2150), .Q(\registers[8][1] )
         );
  DLH_X1 \registers_reg[8][0]  ( .G(n1991), .D(n2153), .Q(\registers[8][0] )
         );
  DLH_X1 \registers_reg[9][31]  ( .G(n1994), .D(n2060), .Q(\registers[9][31] )
         );
  DLH_X1 \registers_reg[9][30]  ( .G(n1994), .D(n2063), .Q(\registers[9][30] )
         );
  DLH_X1 \registers_reg[9][29]  ( .G(n1994), .D(n2066), .Q(\registers[9][29] )
         );
  DLH_X1 \registers_reg[9][28]  ( .G(n1994), .D(n2069), .Q(\registers[9][28] )
         );
  DLH_X1 \registers_reg[9][27]  ( .G(n1994), .D(n2072), .Q(\registers[9][27] )
         );
  DLH_X1 \registers_reg[9][26]  ( .G(n1994), .D(n2075), .Q(\registers[9][26] )
         );
  DLH_X1 \registers_reg[9][25]  ( .G(n1994), .D(n2078), .Q(\registers[9][25] )
         );
  DLH_X1 \registers_reg[9][24]  ( .G(n1993), .D(n2081), .Q(\registers[9][24] )
         );
  DLH_X1 \registers_reg[9][23]  ( .G(n1993), .D(n2084), .Q(\registers[9][23] )
         );
  DLH_X1 \registers_reg[9][22]  ( .G(n1993), .D(n2087), .Q(\registers[9][22] )
         );
  DLH_X1 \registers_reg[9][21]  ( .G(n1993), .D(n2090), .Q(\registers[9][21] )
         );
  DLH_X1 \registers_reg[9][20]  ( .G(n1994), .D(n2093), .Q(\registers[9][20] )
         );
  DLH_X1 \registers_reg[9][19]  ( .G(n1993), .D(n2096), .Q(\registers[9][19] )
         );
  DLH_X1 \registers_reg[9][18]  ( .G(n1993), .D(n2099), .Q(\registers[9][18] )
         );
  DLH_X1 \registers_reg[9][17]  ( .G(n1994), .D(n2102), .Q(\registers[9][17] )
         );
  DLH_X1 \registers_reg[9][16]  ( .G(n1993), .D(n2105), .Q(\registers[9][16] )
         );
  DLH_X1 \registers_reg[9][15]  ( .G(n1993), .D(n2108), .Q(\registers[9][15] )
         );
  DLH_X1 \registers_reg[9][14]  ( .G(n1993), .D(n2111), .Q(\registers[9][14] )
         );
  DLH_X1 \registers_reg[9][13]  ( .G(n1992), .D(n2114), .Q(\registers[9][13] )
         );
  DLH_X1 \registers_reg[9][12]  ( .G(n1993), .D(n2117), .Q(\registers[9][12] )
         );
  DLH_X1 \registers_reg[9][11]  ( .G(n1992), .D(n2120), .Q(\registers[9][11] )
         );
  DLH_X1 \registers_reg[9][10]  ( .G(n1992), .D(n2123), .Q(\registers[9][10] )
         );
  DLH_X1 \registers_reg[9][9]  ( .G(n1992), .D(n2126), .Q(\registers[9][9] )
         );
  DLH_X1 \registers_reg[9][8]  ( .G(n1992), .D(n2129), .Q(\registers[9][8] )
         );
  DLH_X1 \registers_reg[9][7]  ( .G(n1992), .D(n2132), .Q(\registers[9][7] )
         );
  DLH_X1 \registers_reg[9][6]  ( .G(n1992), .D(n2135), .Q(\registers[9][6] )
         );
  DLH_X1 \registers_reg[9][5]  ( .G(n1992), .D(n2138), .Q(\registers[9][5] )
         );
  DLH_X1 \registers_reg[9][4]  ( .G(n1992), .D(n2141), .Q(\registers[9][4] )
         );
  DLH_X1 \registers_reg[9][3]  ( .G(n1992), .D(n2144), .Q(\registers[9][3] )
         );
  DLH_X1 \registers_reg[9][2]  ( .G(n1992), .D(n2147), .Q(\registers[9][2] )
         );
  DLH_X1 \registers_reg[9][1]  ( .G(n1993), .D(n2150), .Q(\registers[9][1] )
         );
  DLH_X1 \registers_reg[9][0]  ( .G(n1994), .D(n2153), .Q(\registers[9][0] )
         );
  DLH_X1 \registers_reg[10][31]  ( .G(n1997), .D(n2059), .Q(
        \registers[10][31] ) );
  DLH_X1 \registers_reg[10][30]  ( .G(n1997), .D(n2062), .Q(
        \registers[10][30] ) );
  DLH_X1 \registers_reg[10][29]  ( .G(n1997), .D(n2065), .Q(
        \registers[10][29] ) );
  DLH_X1 \registers_reg[10][28]  ( .G(n1997), .D(n2068), .Q(
        \registers[10][28] ) );
  DLH_X1 \registers_reg[10][27]  ( .G(n1997), .D(n2071), .Q(
        \registers[10][27] ) );
  DLH_X1 \registers_reg[10][26]  ( .G(n1997), .D(n2074), .Q(
        \registers[10][26] ) );
  DLH_X1 \registers_reg[10][25]  ( .G(n1997), .D(n2077), .Q(
        \registers[10][25] ) );
  DLH_X1 \registers_reg[10][24]  ( .G(n1996), .D(n2080), .Q(
        \registers[10][24] ) );
  DLH_X1 \registers_reg[10][23]  ( .G(n1996), .D(n2083), .Q(
        \registers[10][23] ) );
  DLH_X1 \registers_reg[10][22]  ( .G(n1996), .D(n2086), .Q(
        \registers[10][22] ) );
  DLH_X1 \registers_reg[10][21]  ( .G(n1996), .D(n2089), .Q(
        \registers[10][21] ) );
  DLH_X1 \registers_reg[10][20]  ( .G(n1997), .D(n2092), .Q(
        \registers[10][20] ) );
  DLH_X1 \registers_reg[10][19]  ( .G(n1996), .D(n2095), .Q(
        \registers[10][19] ) );
  DLH_X1 \registers_reg[10][18]  ( .G(n1996), .D(n2098), .Q(
        \registers[10][18] ) );
  DLH_X1 \registers_reg[10][17]  ( .G(n1997), .D(n2101), .Q(
        \registers[10][17] ) );
  DLH_X1 \registers_reg[10][16]  ( .G(n1996), .D(n2104), .Q(
        \registers[10][16] ) );
  DLH_X1 \registers_reg[10][15]  ( .G(n1996), .D(n2107), .Q(
        \registers[10][15] ) );
  DLH_X1 \registers_reg[10][14]  ( .G(n1996), .D(n2110), .Q(
        \registers[10][14] ) );
  DLH_X1 \registers_reg[10][13]  ( .G(n1995), .D(n2113), .Q(
        \registers[10][13] ) );
  DLH_X1 \registers_reg[10][12]  ( .G(n1996), .D(n2116), .Q(
        \registers[10][12] ) );
  DLH_X1 \registers_reg[10][11]  ( .G(n1995), .D(n2119), .Q(
        \registers[10][11] ) );
  DLH_X1 \registers_reg[10][10]  ( .G(n1995), .D(n2122), .Q(
        \registers[10][10] ) );
  DLH_X1 \registers_reg[10][9]  ( .G(n1995), .D(n2125), .Q(\registers[10][9] )
         );
  DLH_X1 \registers_reg[10][8]  ( .G(n1995), .D(n2128), .Q(\registers[10][8] )
         );
  DLH_X1 \registers_reg[10][7]  ( .G(n1995), .D(n2131), .Q(\registers[10][7] )
         );
  DLH_X1 \registers_reg[10][6]  ( .G(n1995), .D(n2134), .Q(\registers[10][6] )
         );
  DLH_X1 \registers_reg[10][5]  ( .G(n1995), .D(n2137), .Q(\registers[10][5] )
         );
  DLH_X1 \registers_reg[10][4]  ( .G(n1995), .D(n2140), .Q(\registers[10][4] )
         );
  DLH_X1 \registers_reg[10][3]  ( .G(n1995), .D(n2143), .Q(\registers[10][3] )
         );
  DLH_X1 \registers_reg[10][2]  ( .G(n1995), .D(n2146), .Q(\registers[10][2] )
         );
  DLH_X1 \registers_reg[10][1]  ( .G(n1996), .D(n2149), .Q(\registers[10][1] )
         );
  DLH_X1 \registers_reg[10][0]  ( .G(n1997), .D(n2152), .Q(\registers[10][0] )
         );
  DLH_X1 \registers_reg[11][31]  ( .G(n2000), .D(n2059), .Q(
        \registers[11][31] ) );
  DLH_X1 \registers_reg[11][30]  ( .G(n2000), .D(n2062), .Q(
        \registers[11][30] ) );
  DLH_X1 \registers_reg[11][29]  ( .G(n2000), .D(n2065), .Q(
        \registers[11][29] ) );
  DLH_X1 \registers_reg[11][28]  ( .G(n2000), .D(n2068), .Q(
        \registers[11][28] ) );
  DLH_X1 \registers_reg[11][27]  ( .G(n2000), .D(n2071), .Q(
        \registers[11][27] ) );
  DLH_X1 \registers_reg[11][26]  ( .G(n2000), .D(n2074), .Q(
        \registers[11][26] ) );
  DLH_X1 \registers_reg[11][25]  ( .G(n2000), .D(n2077), .Q(
        \registers[11][25] ) );
  DLH_X1 \registers_reg[11][24]  ( .G(n1999), .D(n2080), .Q(
        \registers[11][24] ) );
  DLH_X1 \registers_reg[11][23]  ( .G(n1999), .D(n2083), .Q(
        \registers[11][23] ) );
  DLH_X1 \registers_reg[11][22]  ( .G(n1999), .D(n2086), .Q(
        \registers[11][22] ) );
  DLH_X1 \registers_reg[11][21]  ( .G(n1999), .D(n2089), .Q(
        \registers[11][21] ) );
  DLH_X1 \registers_reg[11][20]  ( .G(n2000), .D(n2092), .Q(
        \registers[11][20] ) );
  DLH_X1 \registers_reg[11][19]  ( .G(n1999), .D(n2095), .Q(
        \registers[11][19] ) );
  DLH_X1 \registers_reg[11][18]  ( .G(n1999), .D(n2098), .Q(
        \registers[11][18] ) );
  DLH_X1 \registers_reg[11][17]  ( .G(n2000), .D(n2101), .Q(
        \registers[11][17] ) );
  DLH_X1 \registers_reg[11][16]  ( .G(n1999), .D(n2104), .Q(
        \registers[11][16] ) );
  DLH_X1 \registers_reg[11][15]  ( .G(n1999), .D(n2107), .Q(
        \registers[11][15] ) );
  DLH_X1 \registers_reg[11][14]  ( .G(n1999), .D(n2110), .Q(
        \registers[11][14] ) );
  DLH_X1 \registers_reg[11][13]  ( .G(n1998), .D(n2113), .Q(
        \registers[11][13] ) );
  DLH_X1 \registers_reg[11][12]  ( .G(n1999), .D(n2116), .Q(
        \registers[11][12] ) );
  DLH_X1 \registers_reg[11][11]  ( .G(n1998), .D(n2119), .Q(
        \registers[11][11] ) );
  DLH_X1 \registers_reg[11][10]  ( .G(n1998), .D(n2122), .Q(
        \registers[11][10] ) );
  DLH_X1 \registers_reg[11][9]  ( .G(n1998), .D(n2125), .Q(\registers[11][9] )
         );
  DLH_X1 \registers_reg[11][8]  ( .G(n1998), .D(n2128), .Q(\registers[11][8] )
         );
  DLH_X1 \registers_reg[11][7]  ( .G(n1998), .D(n2131), .Q(\registers[11][7] )
         );
  DLH_X1 \registers_reg[11][6]  ( .G(n1998), .D(n2134), .Q(\registers[11][6] )
         );
  DLH_X1 \registers_reg[11][5]  ( .G(n1998), .D(n2137), .Q(\registers[11][5] )
         );
  DLH_X1 \registers_reg[11][4]  ( .G(n1998), .D(n2140), .Q(\registers[11][4] )
         );
  DLH_X1 \registers_reg[11][3]  ( .G(n1998), .D(n2143), .Q(\registers[11][3] )
         );
  DLH_X1 \registers_reg[11][2]  ( .G(n1998), .D(n2146), .Q(\registers[11][2] )
         );
  DLH_X1 \registers_reg[11][1]  ( .G(n1999), .D(n2149), .Q(\registers[11][1] )
         );
  DLH_X1 \registers_reg[11][0]  ( .G(n2000), .D(n2152), .Q(\registers[11][0] )
         );
  DLH_X1 \registers_reg[12][31]  ( .G(n2001), .D(n2059), .Q(
        \registers[12][31] ) );
  DLH_X1 \registers_reg[12][30]  ( .G(n2001), .D(n2062), .Q(
        \registers[12][30] ) );
  DLH_X1 \registers_reg[12][29]  ( .G(n2001), .D(n2065), .Q(
        \registers[12][29] ) );
  DLH_X1 \registers_reg[12][28]  ( .G(n2001), .D(n2068), .Q(
        \registers[12][28] ) );
  DLH_X1 \registers_reg[12][27]  ( .G(n2001), .D(n2071), .Q(
        \registers[12][27] ) );
  DLH_X1 \registers_reg[12][26]  ( .G(n2001), .D(n2074), .Q(
        \registers[12][26] ) );
  DLH_X1 \registers_reg[12][25]  ( .G(n2001), .D(n2077), .Q(
        \registers[12][25] ) );
  DLH_X1 \registers_reg[12][24]  ( .G(n2002), .D(n2080), .Q(
        \registers[12][24] ) );
  DLH_X1 \registers_reg[12][23]  ( .G(n2002), .D(n2083), .Q(
        \registers[12][23] ) );
  DLH_X1 \registers_reg[12][22]  ( .G(n2002), .D(n2086), .Q(
        \registers[12][22] ) );
  DLH_X1 \registers_reg[12][21]  ( .G(n2002), .D(n2089), .Q(
        \registers[12][21] ) );
  DLH_X1 \registers_reg[12][20]  ( .G(n2001), .D(n2092), .Q(
        \registers[12][20] ) );
  DLH_X1 \registers_reg[12][19]  ( .G(n2002), .D(n2095), .Q(
        \registers[12][19] ) );
  DLH_X1 \registers_reg[12][18]  ( .G(n2002), .D(n2098), .Q(
        \registers[12][18] ) );
  DLH_X1 \registers_reg[12][17]  ( .G(n2001), .D(n2101), .Q(
        \registers[12][17] ) );
  DLH_X1 \registers_reg[12][16]  ( .G(n2002), .D(n2104), .Q(
        \registers[12][16] ) );
  DLH_X1 \registers_reg[12][15]  ( .G(n2002), .D(n2107), .Q(
        \registers[12][15] ) );
  DLH_X1 \registers_reg[12][14]  ( .G(n2002), .D(n2110), .Q(
        \registers[12][14] ) );
  DLH_X1 \registers_reg[12][13]  ( .G(n2002), .D(n2113), .Q(
        \registers[12][13] ) );
  DLH_X1 \registers_reg[12][12]  ( .G(n2002), .D(n2116), .Q(
        \registers[12][12] ) );
  DLH_X1 \registers_reg[12][11]  ( .G(n2003), .D(n2119), .Q(
        \registers[12][11] ) );
  DLH_X1 \registers_reg[12][10]  ( .G(n2003), .D(n2122), .Q(
        \registers[12][10] ) );
  DLH_X1 \registers_reg[12][9]  ( .G(n2003), .D(n2125), .Q(\registers[12][9] )
         );
  DLH_X1 \registers_reg[12][8]  ( .G(n2003), .D(n2128), .Q(\registers[12][8] )
         );
  DLH_X1 \registers_reg[12][7]  ( .G(n2003), .D(n2131), .Q(\registers[12][7] )
         );
  DLH_X1 \registers_reg[12][6]  ( .G(n2003), .D(n2134), .Q(\registers[12][6] )
         );
  DLH_X1 \registers_reg[12][5]  ( .G(n2003), .D(n2137), .Q(\registers[12][5] )
         );
  DLH_X1 \registers_reg[12][4]  ( .G(n2003), .D(n2140), .Q(\registers[12][4] )
         );
  DLH_X1 \registers_reg[12][3]  ( .G(n2003), .D(n2143), .Q(\registers[12][3] )
         );
  DLH_X1 \registers_reg[12][2]  ( .G(n2003), .D(n2146), .Q(\registers[12][2] )
         );
  DLH_X1 \registers_reg[12][1]  ( .G(n2001), .D(n2149), .Q(\registers[12][1] )
         );
  DLH_X1 \registers_reg[12][0]  ( .G(n2001), .D(n2152), .Q(\registers[12][0] )
         );
  DLH_X1 \registers_reg[13][31]  ( .G(n2004), .D(n2059), .Q(
        \registers[13][31] ) );
  DLH_X1 \registers_reg[13][30]  ( .G(n2004), .D(n2062), .Q(
        \registers[13][30] ) );
  DLH_X1 \registers_reg[13][29]  ( .G(n2004), .D(n2065), .Q(
        \registers[13][29] ) );
  DLH_X1 \registers_reg[13][28]  ( .G(n2004), .D(n2068), .Q(
        \registers[13][28] ) );
  DLH_X1 \registers_reg[13][27]  ( .G(n2004), .D(n2071), .Q(
        \registers[13][27] ) );
  DLH_X1 \registers_reg[13][26]  ( .G(n2004), .D(n2074), .Q(
        \registers[13][26] ) );
  DLH_X1 \registers_reg[13][25]  ( .G(n2004), .D(n2077), .Q(
        \registers[13][25] ) );
  DLH_X1 \registers_reg[13][24]  ( .G(n2005), .D(n2080), .Q(
        \registers[13][24] ) );
  DLH_X1 \registers_reg[13][23]  ( .G(n2005), .D(n2083), .Q(
        \registers[13][23] ) );
  DLH_X1 \registers_reg[13][22]  ( .G(n2005), .D(n2086), .Q(
        \registers[13][22] ) );
  DLH_X1 \registers_reg[13][21]  ( .G(n2005), .D(n2089), .Q(
        \registers[13][21] ) );
  DLH_X1 \registers_reg[13][20]  ( .G(n2004), .D(n2092), .Q(
        \registers[13][20] ) );
  DLH_X1 \registers_reg[13][19]  ( .G(n2005), .D(n2095), .Q(
        \registers[13][19] ) );
  DLH_X1 \registers_reg[13][18]  ( .G(n2005), .D(n2098), .Q(
        \registers[13][18] ) );
  DLH_X1 \registers_reg[13][17]  ( .G(n2004), .D(n2101), .Q(
        \registers[13][17] ) );
  DLH_X1 \registers_reg[13][16]  ( .G(n2005), .D(n2104), .Q(
        \registers[13][16] ) );
  DLH_X1 \registers_reg[13][15]  ( .G(n2005), .D(n2107), .Q(
        \registers[13][15] ) );
  DLH_X1 \registers_reg[13][14]  ( .G(n2005), .D(n2110), .Q(
        \registers[13][14] ) );
  DLH_X1 \registers_reg[13][13]  ( .G(n2005), .D(n2113), .Q(
        \registers[13][13] ) );
  DLH_X1 \registers_reg[13][12]  ( .G(n2005), .D(n2116), .Q(
        \registers[13][12] ) );
  DLH_X1 \registers_reg[13][11]  ( .G(n2006), .D(n2119), .Q(
        \registers[13][11] ) );
  DLH_X1 \registers_reg[13][10]  ( .G(n2006), .D(n2122), .Q(
        \registers[13][10] ) );
  DLH_X1 \registers_reg[13][9]  ( .G(n2006), .D(n2125), .Q(\registers[13][9] )
         );
  DLH_X1 \registers_reg[13][8]  ( .G(n2006), .D(n2128), .Q(\registers[13][8] )
         );
  DLH_X1 \registers_reg[13][7]  ( .G(n2006), .D(n2131), .Q(\registers[13][7] )
         );
  DLH_X1 \registers_reg[13][6]  ( .G(n2006), .D(n2134), .Q(\registers[13][6] )
         );
  DLH_X1 \registers_reg[13][5]  ( .G(n2006), .D(n2137), .Q(\registers[13][5] )
         );
  DLH_X1 \registers_reg[13][4]  ( .G(n2006), .D(n2140), .Q(\registers[13][4] )
         );
  DLH_X1 \registers_reg[13][3]  ( .G(n2006), .D(n2143), .Q(\registers[13][3] )
         );
  DLH_X1 \registers_reg[13][2]  ( .G(n2006), .D(n2146), .Q(\registers[13][2] )
         );
  DLH_X1 \registers_reg[13][1]  ( .G(n2004), .D(n2149), .Q(\registers[13][1] )
         );
  DLH_X1 \registers_reg[13][0]  ( .G(n2004), .D(n2152), .Q(\registers[13][0] )
         );
  DLH_X1 \registers_reg[14][31]  ( .G(n2007), .D(n2059), .Q(
        \registers[14][31] ) );
  DLH_X1 \registers_reg[14][30]  ( .G(n2007), .D(n2062), .Q(
        \registers[14][30] ) );
  DLH_X1 \registers_reg[14][29]  ( .G(n2007), .D(n2065), .Q(
        \registers[14][29] ) );
  DLH_X1 \registers_reg[14][28]  ( .G(n2007), .D(n2068), .Q(
        \registers[14][28] ) );
  DLH_X1 \registers_reg[14][27]  ( .G(n2007), .D(n2071), .Q(
        \registers[14][27] ) );
  DLH_X1 \registers_reg[14][26]  ( .G(n2007), .D(n2074), .Q(
        \registers[14][26] ) );
  DLH_X1 \registers_reg[14][25]  ( .G(n2007), .D(n2077), .Q(
        \registers[14][25] ) );
  DLH_X1 \registers_reg[14][24]  ( .G(n2008), .D(n2080), .Q(
        \registers[14][24] ) );
  DLH_X1 \registers_reg[14][23]  ( .G(n2008), .D(n2083), .Q(
        \registers[14][23] ) );
  DLH_X1 \registers_reg[14][22]  ( .G(n2008), .D(n2086), .Q(
        \registers[14][22] ) );
  DLH_X1 \registers_reg[14][21]  ( .G(n2008), .D(n2089), .Q(
        \registers[14][21] ) );
  DLH_X1 \registers_reg[14][20]  ( .G(n2007), .D(n2092), .Q(
        \registers[14][20] ) );
  DLH_X1 \registers_reg[14][19]  ( .G(n2008), .D(n2095), .Q(
        \registers[14][19] ) );
  DLH_X1 \registers_reg[14][18]  ( .G(n2008), .D(n2098), .Q(
        \registers[14][18] ) );
  DLH_X1 \registers_reg[14][17]  ( .G(n2007), .D(n2101), .Q(
        \registers[14][17] ) );
  DLH_X1 \registers_reg[14][16]  ( .G(n2008), .D(n2104), .Q(
        \registers[14][16] ) );
  DLH_X1 \registers_reg[14][15]  ( .G(n2008), .D(n2107), .Q(
        \registers[14][15] ) );
  DLH_X1 \registers_reg[14][14]  ( .G(n2008), .D(n2110), .Q(
        \registers[14][14] ) );
  DLH_X1 \registers_reg[14][13]  ( .G(n2008), .D(n2113), .Q(
        \registers[14][13] ) );
  DLH_X1 \registers_reg[14][12]  ( .G(n2008), .D(n2116), .Q(
        \registers[14][12] ) );
  DLH_X1 \registers_reg[14][11]  ( .G(n2009), .D(n2119), .Q(
        \registers[14][11] ) );
  DLH_X1 \registers_reg[14][10]  ( .G(n2009), .D(n2122), .Q(
        \registers[14][10] ) );
  DLH_X1 \registers_reg[14][9]  ( .G(n2009), .D(n2125), .Q(\registers[14][9] )
         );
  DLH_X1 \registers_reg[14][8]  ( .G(n2009), .D(n2128), .Q(\registers[14][8] )
         );
  DLH_X1 \registers_reg[14][7]  ( .G(n2009), .D(n2131), .Q(\registers[14][7] )
         );
  DLH_X1 \registers_reg[14][6]  ( .G(n2009), .D(n2134), .Q(\registers[14][6] )
         );
  DLH_X1 \registers_reg[14][5]  ( .G(n2009), .D(n2137), .Q(\registers[14][5] )
         );
  DLH_X1 \registers_reg[14][4]  ( .G(n2009), .D(n2140), .Q(\registers[14][4] )
         );
  DLH_X1 \registers_reg[14][3]  ( .G(n2009), .D(n2143), .Q(\registers[14][3] )
         );
  DLH_X1 \registers_reg[14][2]  ( .G(n2009), .D(n2146), .Q(\registers[14][2] )
         );
  DLH_X1 \registers_reg[14][1]  ( .G(n2007), .D(n2149), .Q(\registers[14][1] )
         );
  DLH_X1 \registers_reg[14][0]  ( .G(n2007), .D(n2152), .Q(\registers[14][0] )
         );
  DLH_X1 \registers_reg[15][31]  ( .G(n2010), .D(n2059), .Q(
        \registers[15][31] ) );
  DLH_X1 \registers_reg[15][30]  ( .G(n2010), .D(n2062), .Q(
        \registers[15][30] ) );
  DLH_X1 \registers_reg[15][29]  ( .G(n2010), .D(n2065), .Q(
        \registers[15][29] ) );
  DLH_X1 \registers_reg[15][28]  ( .G(n2010), .D(n2068), .Q(
        \registers[15][28] ) );
  DLH_X1 \registers_reg[15][27]  ( .G(n2010), .D(n2071), .Q(
        \registers[15][27] ) );
  DLH_X1 \registers_reg[15][26]  ( .G(n2010), .D(n2074), .Q(
        \registers[15][26] ) );
  DLH_X1 \registers_reg[15][25]  ( .G(n2010), .D(n2077), .Q(
        \registers[15][25] ) );
  DLH_X1 \registers_reg[15][24]  ( .G(n2011), .D(n2080), .Q(
        \registers[15][24] ) );
  DLH_X1 \registers_reg[15][23]  ( .G(n2011), .D(n2083), .Q(
        \registers[15][23] ) );
  DLH_X1 \registers_reg[15][22]  ( .G(n2011), .D(n2086), .Q(
        \registers[15][22] ) );
  DLH_X1 \registers_reg[15][21]  ( .G(n2011), .D(n2089), .Q(
        \registers[15][21] ) );
  DLH_X1 \registers_reg[15][20]  ( .G(n2010), .D(n2092), .Q(
        \registers[15][20] ) );
  DLH_X1 \registers_reg[15][19]  ( .G(n2011), .D(n2095), .Q(
        \registers[15][19] ) );
  DLH_X1 \registers_reg[15][18]  ( .G(n2011), .D(n2098), .Q(
        \registers[15][18] ) );
  DLH_X1 \registers_reg[15][17]  ( .G(n2010), .D(n2101), .Q(
        \registers[15][17] ) );
  DLH_X1 \registers_reg[15][16]  ( .G(n2011), .D(n2104), .Q(
        \registers[15][16] ) );
  DLH_X1 \registers_reg[15][15]  ( .G(n2011), .D(n2107), .Q(
        \registers[15][15] ) );
  DLH_X1 \registers_reg[15][14]  ( .G(n2011), .D(n2110), .Q(
        \registers[15][14] ) );
  DLH_X1 \registers_reg[15][13]  ( .G(n2011), .D(n2113), .Q(
        \registers[15][13] ) );
  DLH_X1 \registers_reg[15][12]  ( .G(n2011), .D(n2116), .Q(
        \registers[15][12] ) );
  DLH_X1 \registers_reg[15][11]  ( .G(n2012), .D(n2119), .Q(
        \registers[15][11] ) );
  DLH_X1 \registers_reg[15][10]  ( .G(n2012), .D(n2122), .Q(
        \registers[15][10] ) );
  DLH_X1 \registers_reg[15][9]  ( .G(n2012), .D(n2125), .Q(\registers[15][9] )
         );
  DLH_X1 \registers_reg[15][8]  ( .G(n2012), .D(n2128), .Q(\registers[15][8] )
         );
  DLH_X1 \registers_reg[15][7]  ( .G(n2012), .D(n2131), .Q(\registers[15][7] )
         );
  DLH_X1 \registers_reg[15][6]  ( .G(n2012), .D(n2134), .Q(\registers[15][6] )
         );
  DLH_X1 \registers_reg[15][5]  ( .G(n2012), .D(n2137), .Q(\registers[15][5] )
         );
  DLH_X1 \registers_reg[15][4]  ( .G(n2012), .D(n2140), .Q(\registers[15][4] )
         );
  DLH_X1 \registers_reg[15][3]  ( .G(n2012), .D(n2143), .Q(\registers[15][3] )
         );
  DLH_X1 \registers_reg[15][2]  ( .G(n2012), .D(n2146), .Q(\registers[15][2] )
         );
  DLH_X1 \registers_reg[15][1]  ( .G(n2010), .D(n2149), .Q(\registers[15][1] )
         );
  DLH_X1 \registers_reg[15][0]  ( .G(n2010), .D(n2152), .Q(\registers[15][0] )
         );
  DLH_X1 \registers_reg[16][31]  ( .G(n2013), .D(n2059), .Q(
        \registers[16][31] ) );
  DLH_X1 \registers_reg[16][30]  ( .G(n2013), .D(n2062), .Q(
        \registers[16][30] ) );
  DLH_X1 \registers_reg[16][29]  ( .G(n2013), .D(n2065), .Q(
        \registers[16][29] ) );
  DLH_X1 \registers_reg[16][28]  ( .G(n2013), .D(n2068), .Q(
        \registers[16][28] ) );
  DLH_X1 \registers_reg[16][27]  ( .G(n2013), .D(n2071), .Q(
        \registers[16][27] ) );
  DLH_X1 \registers_reg[16][26]  ( .G(n2013), .D(n2074), .Q(
        \registers[16][26] ) );
  DLH_X1 \registers_reg[16][25]  ( .G(n2013), .D(n2077), .Q(
        \registers[16][25] ) );
  DLH_X1 \registers_reg[16][24]  ( .G(n2014), .D(n2080), .Q(
        \registers[16][24] ) );
  DLH_X1 \registers_reg[16][23]  ( .G(n2014), .D(n2083), .Q(
        \registers[16][23] ) );
  DLH_X1 \registers_reg[16][22]  ( .G(n2014), .D(n2086), .Q(
        \registers[16][22] ) );
  DLH_X1 \registers_reg[16][21]  ( .G(n2014), .D(n2089), .Q(
        \registers[16][21] ) );
  DLH_X1 \registers_reg[16][20]  ( .G(n2013), .D(n2092), .Q(
        \registers[16][20] ) );
  DLH_X1 \registers_reg[16][19]  ( .G(n2014), .D(n2095), .Q(
        \registers[16][19] ) );
  DLH_X1 \registers_reg[16][18]  ( .G(n2014), .D(n2098), .Q(
        \registers[16][18] ) );
  DLH_X1 \registers_reg[16][17]  ( .G(n2013), .D(n2101), .Q(
        \registers[16][17] ) );
  DLH_X1 \registers_reg[16][16]  ( .G(n2014), .D(n2104), .Q(
        \registers[16][16] ) );
  DLH_X1 \registers_reg[16][15]  ( .G(n2014), .D(n2107), .Q(
        \registers[16][15] ) );
  DLH_X1 \registers_reg[16][14]  ( .G(n2014), .D(n2110), .Q(
        \registers[16][14] ) );
  DLH_X1 \registers_reg[16][13]  ( .G(n2014), .D(n2113), .Q(
        \registers[16][13] ) );
  DLH_X1 \registers_reg[16][12]  ( .G(n2014), .D(n2116), .Q(
        \registers[16][12] ) );
  DLH_X1 \registers_reg[16][11]  ( .G(n2015), .D(n2119), .Q(
        \registers[16][11] ) );
  DLH_X1 \registers_reg[16][10]  ( .G(n2015), .D(n2122), .Q(
        \registers[16][10] ) );
  DLH_X1 \registers_reg[16][9]  ( .G(n2015), .D(n2125), .Q(\registers[16][9] )
         );
  DLH_X1 \registers_reg[16][8]  ( .G(n2015), .D(n2128), .Q(\registers[16][8] )
         );
  DLH_X1 \registers_reg[16][7]  ( .G(n2015), .D(n2131), .Q(\registers[16][7] )
         );
  DLH_X1 \registers_reg[16][6]  ( .G(n2015), .D(n2134), .Q(\registers[16][6] )
         );
  DLH_X1 \registers_reg[16][5]  ( .G(n2015), .D(n2137), .Q(\registers[16][5] )
         );
  DLH_X1 \registers_reg[16][4]  ( .G(n2015), .D(n2140), .Q(\registers[16][4] )
         );
  DLH_X1 \registers_reg[16][3]  ( .G(n2015), .D(n2143), .Q(\registers[16][3] )
         );
  DLH_X1 \registers_reg[16][2]  ( .G(n2015), .D(n2146), .Q(\registers[16][2] )
         );
  DLH_X1 \registers_reg[16][1]  ( .G(n2013), .D(n2149), .Q(\registers[16][1] )
         );
  DLH_X1 \registers_reg[16][0]  ( .G(n2013), .D(n2152), .Q(\registers[16][0] )
         );
  DLH_X1 \registers_reg[17][31]  ( .G(n2016), .D(n2059), .Q(
        \registers[17][31] ) );
  DLH_X1 \registers_reg[17][30]  ( .G(n2016), .D(n2062), .Q(
        \registers[17][30] ) );
  DLH_X1 \registers_reg[17][29]  ( .G(n2016), .D(n2065), .Q(
        \registers[17][29] ) );
  DLH_X1 \registers_reg[17][28]  ( .G(n2016), .D(n2068), .Q(
        \registers[17][28] ) );
  DLH_X1 \registers_reg[17][27]  ( .G(n2016), .D(n2071), .Q(
        \registers[17][27] ) );
  DLH_X1 \registers_reg[17][26]  ( .G(n2016), .D(n2074), .Q(
        \registers[17][26] ) );
  DLH_X1 \registers_reg[17][25]  ( .G(n2016), .D(n2077), .Q(
        \registers[17][25] ) );
  DLH_X1 \registers_reg[17][24]  ( .G(n2017), .D(n2080), .Q(
        \registers[17][24] ) );
  DLH_X1 \registers_reg[17][23]  ( .G(n2017), .D(n2083), .Q(
        \registers[17][23] ) );
  DLH_X1 \registers_reg[17][22]  ( .G(n2017), .D(n2086), .Q(
        \registers[17][22] ) );
  DLH_X1 \registers_reg[17][21]  ( .G(n2017), .D(n2089), .Q(
        \registers[17][21] ) );
  DLH_X1 \registers_reg[17][20]  ( .G(n2016), .D(n2092), .Q(
        \registers[17][20] ) );
  DLH_X1 \registers_reg[17][19]  ( .G(n2017), .D(n2095), .Q(
        \registers[17][19] ) );
  DLH_X1 \registers_reg[17][18]  ( .G(n2017), .D(n2098), .Q(
        \registers[17][18] ) );
  DLH_X1 \registers_reg[17][17]  ( .G(n2016), .D(n2101), .Q(
        \registers[17][17] ) );
  DLH_X1 \registers_reg[17][16]  ( .G(n2017), .D(n2104), .Q(
        \registers[17][16] ) );
  DLH_X1 \registers_reg[17][15]  ( .G(n2017), .D(n2107), .Q(
        \registers[17][15] ) );
  DLH_X1 \registers_reg[17][14]  ( .G(n2017), .D(n2110), .Q(
        \registers[17][14] ) );
  DLH_X1 \registers_reg[17][13]  ( .G(n2017), .D(n2113), .Q(
        \registers[17][13] ) );
  DLH_X1 \registers_reg[17][12]  ( .G(n2017), .D(n2116), .Q(
        \registers[17][12] ) );
  DLH_X1 \registers_reg[17][11]  ( .G(n2018), .D(n2119), .Q(
        \registers[17][11] ) );
  DLH_X1 \registers_reg[17][10]  ( .G(n2018), .D(n2122), .Q(
        \registers[17][10] ) );
  DLH_X1 \registers_reg[17][9]  ( .G(n2018), .D(n2125), .Q(\registers[17][9] )
         );
  DLH_X1 \registers_reg[17][8]  ( .G(n2018), .D(n2128), .Q(\registers[17][8] )
         );
  DLH_X1 \registers_reg[17][7]  ( .G(n2018), .D(n2131), .Q(\registers[17][7] )
         );
  DLH_X1 \registers_reg[17][6]  ( .G(n2018), .D(n2134), .Q(\registers[17][6] )
         );
  DLH_X1 \registers_reg[17][5]  ( .G(n2018), .D(n2137), .Q(\registers[17][5] )
         );
  DLH_X1 \registers_reg[17][4]  ( .G(n2018), .D(n2140), .Q(\registers[17][4] )
         );
  DLH_X1 \registers_reg[17][3]  ( .G(n2018), .D(n2143), .Q(\registers[17][3] )
         );
  DLH_X1 \registers_reg[17][2]  ( .G(n2018), .D(n2146), .Q(\registers[17][2] )
         );
  DLH_X1 \registers_reg[17][1]  ( .G(n2016), .D(n2149), .Q(\registers[17][1] )
         );
  DLH_X1 \registers_reg[17][0]  ( .G(n2016), .D(n2152), .Q(\registers[17][0] )
         );
  DLH_X1 \registers_reg[18][31]  ( .G(n2019), .D(n2059), .Q(
        \registers[18][31] ) );
  DLH_X1 \registers_reg[18][30]  ( .G(n2019), .D(n2062), .Q(
        \registers[18][30] ) );
  DLH_X1 \registers_reg[18][29]  ( .G(n2019), .D(n2065), .Q(
        \registers[18][29] ) );
  DLH_X1 \registers_reg[18][28]  ( .G(n2019), .D(n2068), .Q(
        \registers[18][28] ) );
  DLH_X1 \registers_reg[18][27]  ( .G(n2019), .D(n2071), .Q(
        \registers[18][27] ) );
  DLH_X1 \registers_reg[18][26]  ( .G(n2019), .D(n2074), .Q(
        \registers[18][26] ) );
  DLH_X1 \registers_reg[18][25]  ( .G(n2019), .D(n2077), .Q(
        \registers[18][25] ) );
  DLH_X1 \registers_reg[18][24]  ( .G(n2020), .D(n2080), .Q(
        \registers[18][24] ) );
  DLH_X1 \registers_reg[18][23]  ( .G(n2020), .D(n2083), .Q(
        \registers[18][23] ) );
  DLH_X1 \registers_reg[18][22]  ( .G(n2020), .D(n2086), .Q(
        \registers[18][22] ) );
  DLH_X1 \registers_reg[18][21]  ( .G(n2020), .D(n2089), .Q(
        \registers[18][21] ) );
  DLH_X1 \registers_reg[18][20]  ( .G(n2019), .D(n2092), .Q(
        \registers[18][20] ) );
  DLH_X1 \registers_reg[18][19]  ( .G(n2020), .D(n2095), .Q(
        \registers[18][19] ) );
  DLH_X1 \registers_reg[18][18]  ( .G(n2020), .D(n2098), .Q(
        \registers[18][18] ) );
  DLH_X1 \registers_reg[18][17]  ( .G(n2019), .D(n2101), .Q(
        \registers[18][17] ) );
  DLH_X1 \registers_reg[18][16]  ( .G(n2020), .D(n2104), .Q(
        \registers[18][16] ) );
  DLH_X1 \registers_reg[18][15]  ( .G(n2020), .D(n2107), .Q(
        \registers[18][15] ) );
  DLH_X1 \registers_reg[18][14]  ( .G(n2020), .D(n2110), .Q(
        \registers[18][14] ) );
  DLH_X1 \registers_reg[18][13]  ( .G(n2020), .D(n2113), .Q(
        \registers[18][13] ) );
  DLH_X1 \registers_reg[18][12]  ( .G(n2020), .D(n2116), .Q(
        \registers[18][12] ) );
  DLH_X1 \registers_reg[18][11]  ( .G(n2021), .D(n2119), .Q(
        \registers[18][11] ) );
  DLH_X1 \registers_reg[18][10]  ( .G(n2021), .D(n2122), .Q(
        \registers[18][10] ) );
  DLH_X1 \registers_reg[18][9]  ( .G(n2021), .D(n2125), .Q(\registers[18][9] )
         );
  DLH_X1 \registers_reg[18][8]  ( .G(n2021), .D(n2128), .Q(\registers[18][8] )
         );
  DLH_X1 \registers_reg[18][7]  ( .G(n2021), .D(n2131), .Q(\registers[18][7] )
         );
  DLH_X1 \registers_reg[18][6]  ( .G(n2021), .D(n2134), .Q(\registers[18][6] )
         );
  DLH_X1 \registers_reg[18][5]  ( .G(n2021), .D(n2137), .Q(\registers[18][5] )
         );
  DLH_X1 \registers_reg[18][4]  ( .G(n2021), .D(n2140), .Q(\registers[18][4] )
         );
  DLH_X1 \registers_reg[18][3]  ( .G(n2021), .D(n2143), .Q(\registers[18][3] )
         );
  DLH_X1 \registers_reg[18][2]  ( .G(n2021), .D(n2146), .Q(\registers[18][2] )
         );
  DLH_X1 \registers_reg[18][1]  ( .G(n2019), .D(n2149), .Q(\registers[18][1] )
         );
  DLH_X1 \registers_reg[18][0]  ( .G(n2019), .D(n2152), .Q(\registers[18][0] )
         );
  DLH_X1 \registers_reg[19][31]  ( .G(n2022), .D(n2059), .Q(
        \registers[19][31] ) );
  DLH_X1 \registers_reg[19][30]  ( .G(n2022), .D(n2062), .Q(
        \registers[19][30] ) );
  DLH_X1 \registers_reg[19][29]  ( .G(n2022), .D(n2065), .Q(
        \registers[19][29] ) );
  DLH_X1 \registers_reg[19][28]  ( .G(n2022), .D(n2068), .Q(
        \registers[19][28] ) );
  DLH_X1 \registers_reg[19][27]  ( .G(n2022), .D(n2071), .Q(
        \registers[19][27] ) );
  DLH_X1 \registers_reg[19][26]  ( .G(n2022), .D(n2074), .Q(
        \registers[19][26] ) );
  DLH_X1 \registers_reg[19][25]  ( .G(n2022), .D(n2077), .Q(
        \registers[19][25] ) );
  DLH_X1 \registers_reg[19][24]  ( .G(n2023), .D(n2080), .Q(
        \registers[19][24] ) );
  DLH_X1 \registers_reg[19][23]  ( .G(n2023), .D(n2083), .Q(
        \registers[19][23] ) );
  DLH_X1 \registers_reg[19][22]  ( .G(n2023), .D(n2086), .Q(
        \registers[19][22] ) );
  DLH_X1 \registers_reg[19][21]  ( .G(n2023), .D(n2089), .Q(
        \registers[19][21] ) );
  DLH_X1 \registers_reg[19][20]  ( .G(n2022), .D(n2092), .Q(
        \registers[19][20] ) );
  DLH_X1 \registers_reg[19][19]  ( .G(n2023), .D(n2095), .Q(
        \registers[19][19] ) );
  DLH_X1 \registers_reg[19][18]  ( .G(n2023), .D(n2098), .Q(
        \registers[19][18] ) );
  DLH_X1 \registers_reg[19][17]  ( .G(n2022), .D(n2101), .Q(
        \registers[19][17] ) );
  DLH_X1 \registers_reg[19][16]  ( .G(n2023), .D(n2104), .Q(
        \registers[19][16] ) );
  DLH_X1 \registers_reg[19][15]  ( .G(n2023), .D(n2107), .Q(
        \registers[19][15] ) );
  DLH_X1 \registers_reg[19][14]  ( .G(n2023), .D(n2110), .Q(
        \registers[19][14] ) );
  DLH_X1 \registers_reg[19][13]  ( .G(n2023), .D(n2113), .Q(
        \registers[19][13] ) );
  DLH_X1 \registers_reg[19][12]  ( .G(n2023), .D(n2116), .Q(
        \registers[19][12] ) );
  DLH_X1 \registers_reg[19][11]  ( .G(n2024), .D(n2119), .Q(
        \registers[19][11] ) );
  DLH_X1 \registers_reg[19][10]  ( .G(n2024), .D(n2122), .Q(
        \registers[19][10] ) );
  DLH_X1 \registers_reg[19][9]  ( .G(n2024), .D(n2125), .Q(\registers[19][9] )
         );
  DLH_X1 \registers_reg[19][8]  ( .G(n2024), .D(n2128), .Q(\registers[19][8] )
         );
  DLH_X1 \registers_reg[19][7]  ( .G(n2024), .D(n2131), .Q(\registers[19][7] )
         );
  DLH_X1 \registers_reg[19][6]  ( .G(n2024), .D(n2134), .Q(\registers[19][6] )
         );
  DLH_X1 \registers_reg[19][5]  ( .G(n2024), .D(n2137), .Q(\registers[19][5] )
         );
  DLH_X1 \registers_reg[19][4]  ( .G(n2024), .D(n2140), .Q(\registers[19][4] )
         );
  DLH_X1 \registers_reg[19][3]  ( .G(n2024), .D(n2143), .Q(\registers[19][3] )
         );
  DLH_X1 \registers_reg[19][2]  ( .G(n2024), .D(n2146), .Q(\registers[19][2] )
         );
  DLH_X1 \registers_reg[19][1]  ( .G(n2022), .D(n2149), .Q(\registers[19][1] )
         );
  DLH_X1 \registers_reg[19][0]  ( .G(n2022), .D(n2152), .Q(\registers[19][0] )
         );
  DLH_X1 \registers_reg[20][31]  ( .G(n2025), .D(n2059), .Q(
        \registers[20][31] ) );
  DLH_X1 \registers_reg[20][30]  ( .G(n2025), .D(n2062), .Q(
        \registers[20][30] ) );
  DLH_X1 \registers_reg[20][29]  ( .G(n2025), .D(n2065), .Q(
        \registers[20][29] ) );
  DLH_X1 \registers_reg[20][28]  ( .G(n2025), .D(n2068), .Q(
        \registers[20][28] ) );
  DLH_X1 \registers_reg[20][27]  ( .G(n2025), .D(n2071), .Q(
        \registers[20][27] ) );
  DLH_X1 \registers_reg[20][26]  ( .G(n2025), .D(n2074), .Q(
        \registers[20][26] ) );
  DLH_X1 \registers_reg[20][25]  ( .G(n2025), .D(n2077), .Q(
        \registers[20][25] ) );
  DLH_X1 \registers_reg[20][24]  ( .G(n2026), .D(n2080), .Q(
        \registers[20][24] ) );
  DLH_X1 \registers_reg[20][23]  ( .G(n2026), .D(n2083), .Q(
        \registers[20][23] ) );
  DLH_X1 \registers_reg[20][22]  ( .G(n2026), .D(n2086), .Q(
        \registers[20][22] ) );
  DLH_X1 \registers_reg[20][21]  ( .G(n2026), .D(n2089), .Q(
        \registers[20][21] ) );
  DLH_X1 \registers_reg[20][20]  ( .G(n2025), .D(n2092), .Q(
        \registers[20][20] ) );
  DLH_X1 \registers_reg[20][19]  ( .G(n2026), .D(n2095), .Q(
        \registers[20][19] ) );
  DLH_X1 \registers_reg[20][18]  ( .G(n2026), .D(n2098), .Q(
        \registers[20][18] ) );
  DLH_X1 \registers_reg[20][17]  ( .G(n2025), .D(n2101), .Q(
        \registers[20][17] ) );
  DLH_X1 \registers_reg[20][16]  ( .G(n2026), .D(n2104), .Q(
        \registers[20][16] ) );
  DLH_X1 \registers_reg[20][15]  ( .G(n2026), .D(n2107), .Q(
        \registers[20][15] ) );
  DLH_X1 \registers_reg[20][14]  ( .G(n2026), .D(n2110), .Q(
        \registers[20][14] ) );
  DLH_X1 \registers_reg[20][13]  ( .G(n2026), .D(n2113), .Q(
        \registers[20][13] ) );
  DLH_X1 \registers_reg[20][12]  ( .G(n2026), .D(n2116), .Q(
        \registers[20][12] ) );
  DLH_X1 \registers_reg[20][11]  ( .G(n2027), .D(n2119), .Q(
        \registers[20][11] ) );
  DLH_X1 \registers_reg[20][10]  ( .G(n2027), .D(n2122), .Q(
        \registers[20][10] ) );
  DLH_X1 \registers_reg[20][9]  ( .G(n2027), .D(n2125), .Q(\registers[20][9] )
         );
  DLH_X1 \registers_reg[20][8]  ( .G(n2027), .D(n2128), .Q(\registers[20][8] )
         );
  DLH_X1 \registers_reg[20][7]  ( .G(n2027), .D(n2131), .Q(\registers[20][7] )
         );
  DLH_X1 \registers_reg[20][6]  ( .G(n2027), .D(n2134), .Q(\registers[20][6] )
         );
  DLH_X1 \registers_reg[20][5]  ( .G(n2027), .D(n2137), .Q(\registers[20][5] )
         );
  DLH_X1 \registers_reg[20][4]  ( .G(n2027), .D(n2140), .Q(\registers[20][4] )
         );
  DLH_X1 \registers_reg[20][3]  ( .G(n2027), .D(n2143), .Q(\registers[20][3] )
         );
  DLH_X1 \registers_reg[20][2]  ( .G(n2027), .D(n2146), .Q(\registers[20][2] )
         );
  DLH_X1 \registers_reg[20][1]  ( .G(n2025), .D(n2149), .Q(\registers[20][1] )
         );
  DLH_X1 \registers_reg[20][0]  ( .G(n2025), .D(n2152), .Q(\registers[20][0] )
         );
  DLH_X1 \registers_reg[21][31]  ( .G(n2028), .D(n2058), .Q(
        \registers[21][31] ) );
  DLH_X1 \registers_reg[21][30]  ( .G(n2028), .D(n2061), .Q(
        \registers[21][30] ) );
  DLH_X1 \registers_reg[21][29]  ( .G(n2028), .D(n2064), .Q(
        \registers[21][29] ) );
  DLH_X1 \registers_reg[21][28]  ( .G(n2028), .D(n2067), .Q(
        \registers[21][28] ) );
  DLH_X1 \registers_reg[21][27]  ( .G(n2028), .D(n2070), .Q(
        \registers[21][27] ) );
  DLH_X1 \registers_reg[21][26]  ( .G(n2028), .D(n2073), .Q(
        \registers[21][26] ) );
  DLH_X1 \registers_reg[21][25]  ( .G(n2028), .D(n2076), .Q(
        \registers[21][25] ) );
  DLH_X1 \registers_reg[21][24]  ( .G(n2029), .D(n2079), .Q(
        \registers[21][24] ) );
  DLH_X1 \registers_reg[21][23]  ( .G(n2029), .D(n2082), .Q(
        \registers[21][23] ) );
  DLH_X1 \registers_reg[21][22]  ( .G(n2029), .D(n2085), .Q(
        \registers[21][22] ) );
  DLH_X1 \registers_reg[21][21]  ( .G(n2029), .D(n2088), .Q(
        \registers[21][21] ) );
  DLH_X1 \registers_reg[21][20]  ( .G(n2028), .D(n2091), .Q(
        \registers[21][20] ) );
  DLH_X1 \registers_reg[21][19]  ( .G(n2029), .D(n2094), .Q(
        \registers[21][19] ) );
  DLH_X1 \registers_reg[21][18]  ( .G(n2029), .D(n2097), .Q(
        \registers[21][18] ) );
  DLH_X1 \registers_reg[21][17]  ( .G(n2028), .D(n2100), .Q(
        \registers[21][17] ) );
  DLH_X1 \registers_reg[21][16]  ( .G(n2029), .D(n2103), .Q(
        \registers[21][16] ) );
  DLH_X1 \registers_reg[21][15]  ( .G(n2029), .D(n2106), .Q(
        \registers[21][15] ) );
  DLH_X1 \registers_reg[21][14]  ( .G(n2029), .D(n2109), .Q(
        \registers[21][14] ) );
  DLH_X1 \registers_reg[21][13]  ( .G(n2029), .D(n2112), .Q(
        \registers[21][13] ) );
  DLH_X1 \registers_reg[21][12]  ( .G(n2029), .D(n2115), .Q(
        \registers[21][12] ) );
  DLH_X1 \registers_reg[21][11]  ( .G(n2030), .D(n2118), .Q(
        \registers[21][11] ) );
  DLH_X1 \registers_reg[21][10]  ( .G(n2030), .D(n2121), .Q(
        \registers[21][10] ) );
  DLH_X1 \registers_reg[21][9]  ( .G(n2030), .D(n2124), .Q(\registers[21][9] )
         );
  DLH_X1 \registers_reg[21][8]  ( .G(n2030), .D(n2127), .Q(\registers[21][8] )
         );
  DLH_X1 \registers_reg[21][7]  ( .G(n2030), .D(n2130), .Q(\registers[21][7] )
         );
  DLH_X1 \registers_reg[21][6]  ( .G(n2030), .D(n2133), .Q(\registers[21][6] )
         );
  DLH_X1 \registers_reg[21][5]  ( .G(n2030), .D(n2136), .Q(\registers[21][5] )
         );
  DLH_X1 \registers_reg[21][4]  ( .G(n2030), .D(n2139), .Q(\registers[21][4] )
         );
  DLH_X1 \registers_reg[21][3]  ( .G(n2030), .D(n2142), .Q(\registers[21][3] )
         );
  DLH_X1 \registers_reg[21][2]  ( .G(n2030), .D(n2145), .Q(\registers[21][2] )
         );
  DLH_X1 \registers_reg[21][1]  ( .G(n2028), .D(n2148), .Q(\registers[21][1] )
         );
  DLH_X1 \registers_reg[21][0]  ( .G(n2028), .D(n2151), .Q(\registers[21][0] )
         );
  DLH_X1 \registers_reg[22][31]  ( .G(n2031), .D(n2058), .Q(
        \registers[22][31] ) );
  DLH_X1 \registers_reg[22][30]  ( .G(n2031), .D(n2061), .Q(
        \registers[22][30] ) );
  DLH_X1 \registers_reg[22][29]  ( .G(n2031), .D(n2064), .Q(
        \registers[22][29] ) );
  DLH_X1 \registers_reg[22][28]  ( .G(n2031), .D(n2067), .Q(
        \registers[22][28] ) );
  DLH_X1 \registers_reg[22][27]  ( .G(n2031), .D(n2070), .Q(
        \registers[22][27] ) );
  DLH_X1 \registers_reg[22][26]  ( .G(n2031), .D(n2073), .Q(
        \registers[22][26] ) );
  DLH_X1 \registers_reg[22][25]  ( .G(n2031), .D(n2076), .Q(
        \registers[22][25] ) );
  DLH_X1 \registers_reg[22][24]  ( .G(n2032), .D(n2079), .Q(
        \registers[22][24] ) );
  DLH_X1 \registers_reg[22][23]  ( .G(n2032), .D(n2082), .Q(
        \registers[22][23] ) );
  DLH_X1 \registers_reg[22][22]  ( .G(n2032), .D(n2085), .Q(
        \registers[22][22] ) );
  DLH_X1 \registers_reg[22][21]  ( .G(n2032), .D(n2088), .Q(
        \registers[22][21] ) );
  DLH_X1 \registers_reg[22][20]  ( .G(n2031), .D(n2091), .Q(
        \registers[22][20] ) );
  DLH_X1 \registers_reg[22][19]  ( .G(n2032), .D(n2094), .Q(
        \registers[22][19] ) );
  DLH_X1 \registers_reg[22][18]  ( .G(n2032), .D(n2097), .Q(
        \registers[22][18] ) );
  DLH_X1 \registers_reg[22][17]  ( .G(n2031), .D(n2100), .Q(
        \registers[22][17] ) );
  DLH_X1 \registers_reg[22][16]  ( .G(n2032), .D(n2103), .Q(
        \registers[22][16] ) );
  DLH_X1 \registers_reg[22][15]  ( .G(n2032), .D(n2106), .Q(
        \registers[22][15] ) );
  DLH_X1 \registers_reg[22][14]  ( .G(n2032), .D(n2109), .Q(
        \registers[22][14] ) );
  DLH_X1 \registers_reg[22][13]  ( .G(n2032), .D(n2112), .Q(
        \registers[22][13] ) );
  DLH_X1 \registers_reg[22][12]  ( .G(n2032), .D(n2115), .Q(
        \registers[22][12] ) );
  DLH_X1 \registers_reg[22][11]  ( .G(n2033), .D(n2118), .Q(
        \registers[22][11] ) );
  DLH_X1 \registers_reg[22][10]  ( .G(n2033), .D(n2121), .Q(
        \registers[22][10] ) );
  DLH_X1 \registers_reg[22][9]  ( .G(n2033), .D(n2124), .Q(\registers[22][9] )
         );
  DLH_X1 \registers_reg[22][8]  ( .G(n2033), .D(n2127), .Q(\registers[22][8] )
         );
  DLH_X1 \registers_reg[22][7]  ( .G(n2033), .D(n2130), .Q(\registers[22][7] )
         );
  DLH_X1 \registers_reg[22][6]  ( .G(n2033), .D(n2133), .Q(\registers[22][6] )
         );
  DLH_X1 \registers_reg[22][5]  ( .G(n2033), .D(n2136), .Q(\registers[22][5] )
         );
  DLH_X1 \registers_reg[22][4]  ( .G(n2033), .D(n2139), .Q(\registers[22][4] )
         );
  DLH_X1 \registers_reg[22][3]  ( .G(n2033), .D(n2142), .Q(\registers[22][3] )
         );
  DLH_X1 \registers_reg[22][2]  ( .G(n2033), .D(n2145), .Q(\registers[22][2] )
         );
  DLH_X1 \registers_reg[22][1]  ( .G(n2031), .D(n2148), .Q(\registers[22][1] )
         );
  DLH_X1 \registers_reg[22][0]  ( .G(n2031), .D(n2151), .Q(\registers[22][0] )
         );
  DLH_X1 \registers_reg[23][31]  ( .G(n2034), .D(n2058), .Q(
        \registers[23][31] ) );
  DLH_X1 \registers_reg[23][30]  ( .G(n2034), .D(n2061), .Q(
        \registers[23][30] ) );
  DLH_X1 \registers_reg[23][29]  ( .G(n2034), .D(n2064), .Q(
        \registers[23][29] ) );
  DLH_X1 \registers_reg[23][28]  ( .G(n2034), .D(n2067), .Q(
        \registers[23][28] ) );
  DLH_X1 \registers_reg[23][27]  ( .G(n2034), .D(n2070), .Q(
        \registers[23][27] ) );
  DLH_X1 \registers_reg[23][26]  ( .G(n2034), .D(n2073), .Q(
        \registers[23][26] ) );
  DLH_X1 \registers_reg[23][25]  ( .G(n2034), .D(n2076), .Q(
        \registers[23][25] ) );
  DLH_X1 \registers_reg[23][24]  ( .G(n2035), .D(n2079), .Q(
        \registers[23][24] ) );
  DLH_X1 \registers_reg[23][23]  ( .G(n2035), .D(n2082), .Q(
        \registers[23][23] ) );
  DLH_X1 \registers_reg[23][22]  ( .G(n2035), .D(n2085), .Q(
        \registers[23][22] ) );
  DLH_X1 \registers_reg[23][21]  ( .G(n2035), .D(n2088), .Q(
        \registers[23][21] ) );
  DLH_X1 \registers_reg[23][20]  ( .G(n2034), .D(n2091), .Q(
        \registers[23][20] ) );
  DLH_X1 \registers_reg[23][19]  ( .G(n2035), .D(n2094), .Q(
        \registers[23][19] ) );
  DLH_X1 \registers_reg[23][18]  ( .G(n2035), .D(n2097), .Q(
        \registers[23][18] ) );
  DLH_X1 \registers_reg[23][17]  ( .G(n2034), .D(n2100), .Q(
        \registers[23][17] ) );
  DLH_X1 \registers_reg[23][16]  ( .G(n2035), .D(n2103), .Q(
        \registers[23][16] ) );
  DLH_X1 \registers_reg[23][15]  ( .G(n2035), .D(n2106), .Q(
        \registers[23][15] ) );
  DLH_X1 \registers_reg[23][14]  ( .G(n2035), .D(n2109), .Q(
        \registers[23][14] ) );
  DLH_X1 \registers_reg[23][13]  ( .G(n2035), .D(n2112), .Q(
        \registers[23][13] ) );
  DLH_X1 \registers_reg[23][12]  ( .G(n2035), .D(n2115), .Q(
        \registers[23][12] ) );
  DLH_X1 \registers_reg[23][11]  ( .G(n2036), .D(n2118), .Q(
        \registers[23][11] ) );
  DLH_X1 \registers_reg[23][10]  ( .G(n2036), .D(n2121), .Q(
        \registers[23][10] ) );
  DLH_X1 \registers_reg[23][9]  ( .G(n2036), .D(n2124), .Q(\registers[23][9] )
         );
  DLH_X1 \registers_reg[23][8]  ( .G(n2036), .D(n2127), .Q(\registers[23][8] )
         );
  DLH_X1 \registers_reg[23][7]  ( .G(n2036), .D(n2130), .Q(\registers[23][7] )
         );
  DLH_X1 \registers_reg[23][6]  ( .G(n2036), .D(n2133), .Q(\registers[23][6] )
         );
  DLH_X1 \registers_reg[23][5]  ( .G(n2036), .D(n2136), .Q(\registers[23][5] )
         );
  DLH_X1 \registers_reg[23][4]  ( .G(n2036), .D(n2139), .Q(\registers[23][4] )
         );
  DLH_X1 \registers_reg[23][3]  ( .G(n2036), .D(n2142), .Q(\registers[23][3] )
         );
  DLH_X1 \registers_reg[23][2]  ( .G(n2036), .D(n2145), .Q(\registers[23][2] )
         );
  DLH_X1 \registers_reg[23][1]  ( .G(n2034), .D(n2148), .Q(\registers[23][1] )
         );
  DLH_X1 \registers_reg[23][0]  ( .G(n2034), .D(n2151), .Q(\registers[23][0] )
         );
  DLH_X1 \registers_reg[24][31]  ( .G(n2037), .D(n2058), .Q(
        \registers[24][31] ) );
  DLH_X1 \registers_reg[24][30]  ( .G(n2037), .D(n2061), .Q(
        \registers[24][30] ) );
  DLH_X1 \registers_reg[24][29]  ( .G(n2037), .D(n2064), .Q(
        \registers[24][29] ) );
  DLH_X1 \registers_reg[24][28]  ( .G(n2037), .D(n2067), .Q(
        \registers[24][28] ) );
  DLH_X1 \registers_reg[24][27]  ( .G(n2037), .D(n2070), .Q(
        \registers[24][27] ) );
  DLH_X1 \registers_reg[24][26]  ( .G(n2037), .D(n2073), .Q(
        \registers[24][26] ) );
  DLH_X1 \registers_reg[24][25]  ( .G(n2037), .D(n2076), .Q(
        \registers[24][25] ) );
  DLH_X1 \registers_reg[24][24]  ( .G(n2038), .D(n2079), .Q(
        \registers[24][24] ) );
  DLH_X1 \registers_reg[24][23]  ( .G(n2038), .D(n2082), .Q(
        \registers[24][23] ) );
  DLH_X1 \registers_reg[24][22]  ( .G(n2038), .D(n2085), .Q(
        \registers[24][22] ) );
  DLH_X1 \registers_reg[24][21]  ( .G(n2038), .D(n2088), .Q(
        \registers[24][21] ) );
  DLH_X1 \registers_reg[24][20]  ( .G(n2037), .D(n2091), .Q(
        \registers[24][20] ) );
  DLH_X1 \registers_reg[24][19]  ( .G(n2038), .D(n2094), .Q(
        \registers[24][19] ) );
  DLH_X1 \registers_reg[24][18]  ( .G(n2038), .D(n2097), .Q(
        \registers[24][18] ) );
  DLH_X1 \registers_reg[24][17]  ( .G(n2037), .D(n2100), .Q(
        \registers[24][17] ) );
  DLH_X1 \registers_reg[24][16]  ( .G(n2038), .D(n2103), .Q(
        \registers[24][16] ) );
  DLH_X1 \registers_reg[24][15]  ( .G(n2038), .D(n2106), .Q(
        \registers[24][15] ) );
  DLH_X1 \registers_reg[24][14]  ( .G(n2038), .D(n2109), .Q(
        \registers[24][14] ) );
  DLH_X1 \registers_reg[24][13]  ( .G(n2038), .D(n2112), .Q(
        \registers[24][13] ) );
  DLH_X1 \registers_reg[24][12]  ( .G(n2038), .D(n2115), .Q(
        \registers[24][12] ) );
  DLH_X1 \registers_reg[24][11]  ( .G(n2039), .D(n2118), .Q(
        \registers[24][11] ) );
  DLH_X1 \registers_reg[24][10]  ( .G(n2039), .D(n2121), .Q(
        \registers[24][10] ) );
  DLH_X1 \registers_reg[24][9]  ( .G(n2039), .D(n2124), .Q(\registers[24][9] )
         );
  DLH_X1 \registers_reg[24][8]  ( .G(n2039), .D(n2127), .Q(\registers[24][8] )
         );
  DLH_X1 \registers_reg[24][7]  ( .G(n2039), .D(n2130), .Q(\registers[24][7] )
         );
  DLH_X1 \registers_reg[24][6]  ( .G(n2039), .D(n2133), .Q(\registers[24][6] )
         );
  DLH_X1 \registers_reg[24][5]  ( .G(n2039), .D(n2136), .Q(\registers[24][5] )
         );
  DLH_X1 \registers_reg[24][4]  ( .G(n2039), .D(n2139), .Q(\registers[24][4] )
         );
  DLH_X1 \registers_reg[24][3]  ( .G(n2039), .D(n2142), .Q(\registers[24][3] )
         );
  DLH_X1 \registers_reg[24][2]  ( .G(n2039), .D(n2145), .Q(\registers[24][2] )
         );
  DLH_X1 \registers_reg[24][1]  ( .G(n2037), .D(n2148), .Q(\registers[24][1] )
         );
  DLH_X1 \registers_reg[24][0]  ( .G(n2037), .D(n2151), .Q(\registers[24][0] )
         );
  DLH_X1 \registers_reg[25][31]  ( .G(n2040), .D(n2058), .Q(
        \registers[25][31] ) );
  DLH_X1 \registers_reg[25][30]  ( .G(n2040), .D(n2061), .Q(
        \registers[25][30] ) );
  DLH_X1 \registers_reg[25][29]  ( .G(n2040), .D(n2064), .Q(
        \registers[25][29] ) );
  DLH_X1 \registers_reg[25][28]  ( .G(n2040), .D(n2067), .Q(
        \registers[25][28] ) );
  DLH_X1 \registers_reg[25][27]  ( .G(n2040), .D(n2070), .Q(
        \registers[25][27] ) );
  DLH_X1 \registers_reg[25][26]  ( .G(n2040), .D(n2073), .Q(
        \registers[25][26] ) );
  DLH_X1 \registers_reg[25][25]  ( .G(n2040), .D(n2076), .Q(
        \registers[25][25] ) );
  DLH_X1 \registers_reg[25][24]  ( .G(n2041), .D(n2079), .Q(
        \registers[25][24] ) );
  DLH_X1 \registers_reg[25][23]  ( .G(n2041), .D(n2082), .Q(
        \registers[25][23] ) );
  DLH_X1 \registers_reg[25][22]  ( .G(n2041), .D(n2085), .Q(
        \registers[25][22] ) );
  DLH_X1 \registers_reg[25][21]  ( .G(n2041), .D(n2088), .Q(
        \registers[25][21] ) );
  DLH_X1 \registers_reg[25][20]  ( .G(n2040), .D(n2091), .Q(
        \registers[25][20] ) );
  DLH_X1 \registers_reg[25][19]  ( .G(n2041), .D(n2094), .Q(
        \registers[25][19] ) );
  DLH_X1 \registers_reg[25][18]  ( .G(n2041), .D(n2097), .Q(
        \registers[25][18] ) );
  DLH_X1 \registers_reg[25][17]  ( .G(n2040), .D(n2100), .Q(
        \registers[25][17] ) );
  DLH_X1 \registers_reg[25][16]  ( .G(n2041), .D(n2103), .Q(
        \registers[25][16] ) );
  DLH_X1 \registers_reg[25][15]  ( .G(n2041), .D(n2106), .Q(
        \registers[25][15] ) );
  DLH_X1 \registers_reg[25][14]  ( .G(n2041), .D(n2109), .Q(
        \registers[25][14] ) );
  DLH_X1 \registers_reg[25][13]  ( .G(n2041), .D(n2112), .Q(
        \registers[25][13] ) );
  DLH_X1 \registers_reg[25][12]  ( .G(n2041), .D(n2115), .Q(
        \registers[25][12] ) );
  DLH_X1 \registers_reg[25][11]  ( .G(n2042), .D(n2118), .Q(
        \registers[25][11] ) );
  DLH_X1 \registers_reg[25][10]  ( .G(n2042), .D(n2121), .Q(
        \registers[25][10] ) );
  DLH_X1 \registers_reg[25][9]  ( .G(n2042), .D(n2124), .Q(\registers[25][9] )
         );
  DLH_X1 \registers_reg[25][8]  ( .G(n2042), .D(n2127), .Q(\registers[25][8] )
         );
  DLH_X1 \registers_reg[25][7]  ( .G(n2042), .D(n2130), .Q(\registers[25][7] )
         );
  DLH_X1 \registers_reg[25][6]  ( .G(n2042), .D(n2133), .Q(\registers[25][6] )
         );
  DLH_X1 \registers_reg[25][5]  ( .G(n2042), .D(n2136), .Q(\registers[25][5] )
         );
  DLH_X1 \registers_reg[25][4]  ( .G(n2042), .D(n2139), .Q(\registers[25][4] )
         );
  DLH_X1 \registers_reg[25][3]  ( .G(n2042), .D(n2142), .Q(\registers[25][3] )
         );
  DLH_X1 \registers_reg[25][2]  ( .G(n2042), .D(n2145), .Q(\registers[25][2] )
         );
  DLH_X1 \registers_reg[25][1]  ( .G(n2040), .D(n2148), .Q(\registers[25][1] )
         );
  DLH_X1 \registers_reg[25][0]  ( .G(n2040), .D(n2151), .Q(\registers[25][0] )
         );
  DLH_X1 \registers_reg[26][31]  ( .G(n2043), .D(n2058), .Q(
        \registers[26][31] ) );
  DLH_X1 \registers_reg[26][30]  ( .G(n2043), .D(n2061), .Q(
        \registers[26][30] ) );
  DLH_X1 \registers_reg[26][29]  ( .G(n2043), .D(n2064), .Q(
        \registers[26][29] ) );
  DLH_X1 \registers_reg[26][28]  ( .G(n2043), .D(n2067), .Q(
        \registers[26][28] ) );
  DLH_X1 \registers_reg[26][27]  ( .G(n2043), .D(n2070), .Q(
        \registers[26][27] ) );
  DLH_X1 \registers_reg[26][26]  ( .G(n2043), .D(n2073), .Q(
        \registers[26][26] ) );
  DLH_X1 \registers_reg[26][25]  ( .G(n2043), .D(n2076), .Q(
        \registers[26][25] ) );
  DLH_X1 \registers_reg[26][24]  ( .G(n2044), .D(n2079), .Q(
        \registers[26][24] ) );
  DLH_X1 \registers_reg[26][23]  ( .G(n2044), .D(n2082), .Q(
        \registers[26][23] ) );
  DLH_X1 \registers_reg[26][22]  ( .G(n2044), .D(n2085), .Q(
        \registers[26][22] ) );
  DLH_X1 \registers_reg[26][21]  ( .G(n2044), .D(n2088), .Q(
        \registers[26][21] ) );
  DLH_X1 \registers_reg[26][20]  ( .G(n2043), .D(n2091), .Q(
        \registers[26][20] ) );
  DLH_X1 \registers_reg[26][19]  ( .G(n2044), .D(n2094), .Q(
        \registers[26][19] ) );
  DLH_X1 \registers_reg[26][18]  ( .G(n2044), .D(n2097), .Q(
        \registers[26][18] ) );
  DLH_X1 \registers_reg[26][17]  ( .G(n2043), .D(n2100), .Q(
        \registers[26][17] ) );
  DLH_X1 \registers_reg[26][16]  ( .G(n2044), .D(n2103), .Q(
        \registers[26][16] ) );
  DLH_X1 \registers_reg[26][15]  ( .G(n2044), .D(n2106), .Q(
        \registers[26][15] ) );
  DLH_X1 \registers_reg[26][14]  ( .G(n2044), .D(n2109), .Q(
        \registers[26][14] ) );
  DLH_X1 \registers_reg[26][13]  ( .G(n2044), .D(n2112), .Q(
        \registers[26][13] ) );
  DLH_X1 \registers_reg[26][12]  ( .G(n2044), .D(n2115), .Q(
        \registers[26][12] ) );
  DLH_X1 \registers_reg[26][11]  ( .G(n2045), .D(n2118), .Q(
        \registers[26][11] ) );
  DLH_X1 \registers_reg[26][10]  ( .G(n2045), .D(n2121), .Q(
        \registers[26][10] ) );
  DLH_X1 \registers_reg[26][9]  ( .G(n2045), .D(n2124), .Q(\registers[26][9] )
         );
  DLH_X1 \registers_reg[26][8]  ( .G(n2045), .D(n2127), .Q(\registers[26][8] )
         );
  DLH_X1 \registers_reg[26][7]  ( .G(n2045), .D(n2130), .Q(\registers[26][7] )
         );
  DLH_X1 \registers_reg[26][6]  ( .G(n2045), .D(n2133), .Q(\registers[26][6] )
         );
  DLH_X1 \registers_reg[26][5]  ( .G(n2045), .D(n2136), .Q(\registers[26][5] )
         );
  DLH_X1 \registers_reg[26][4]  ( .G(n2045), .D(n2139), .Q(\registers[26][4] )
         );
  DLH_X1 \registers_reg[26][3]  ( .G(n2045), .D(n2142), .Q(\registers[26][3] )
         );
  DLH_X1 \registers_reg[26][2]  ( .G(n2045), .D(n2145), .Q(\registers[26][2] )
         );
  DLH_X1 \registers_reg[26][1]  ( .G(n2043), .D(n2148), .Q(\registers[26][1] )
         );
  DLH_X1 \registers_reg[26][0]  ( .G(n2043), .D(n2151), .Q(\registers[26][0] )
         );
  DLH_X1 \registers_reg[27][31]  ( .G(n2046), .D(n2058), .Q(
        \registers[27][31] ) );
  DLH_X1 \registers_reg[27][30]  ( .G(n2046), .D(n2061), .Q(
        \registers[27][30] ) );
  DLH_X1 \registers_reg[27][29]  ( .G(n2046), .D(n2064), .Q(
        \registers[27][29] ) );
  DLH_X1 \registers_reg[27][28]  ( .G(n2046), .D(n2067), .Q(
        \registers[27][28] ) );
  DLH_X1 \registers_reg[27][27]  ( .G(n2046), .D(n2070), .Q(
        \registers[27][27] ) );
  DLH_X1 \registers_reg[27][26]  ( .G(n2046), .D(n2073), .Q(
        \registers[27][26] ) );
  DLH_X1 \registers_reg[27][25]  ( .G(n2046), .D(n2076), .Q(
        \registers[27][25] ) );
  DLH_X1 \registers_reg[27][24]  ( .G(n2047), .D(n2079), .Q(
        \registers[27][24] ) );
  DLH_X1 \registers_reg[27][23]  ( .G(n2047), .D(n2082), .Q(
        \registers[27][23] ) );
  DLH_X1 \registers_reg[27][22]  ( .G(n2047), .D(n2085), .Q(
        \registers[27][22] ) );
  DLH_X1 \registers_reg[27][21]  ( .G(n2047), .D(n2088), .Q(
        \registers[27][21] ) );
  DLH_X1 \registers_reg[27][20]  ( .G(n2046), .D(n2091), .Q(
        \registers[27][20] ) );
  DLH_X1 \registers_reg[27][19]  ( .G(n2047), .D(n2094), .Q(
        \registers[27][19] ) );
  DLH_X1 \registers_reg[27][18]  ( .G(n2047), .D(n2097), .Q(
        \registers[27][18] ) );
  DLH_X1 \registers_reg[27][17]  ( .G(n2046), .D(n2100), .Q(
        \registers[27][17] ) );
  DLH_X1 \registers_reg[27][16]  ( .G(n2047), .D(n2103), .Q(
        \registers[27][16] ) );
  DLH_X1 \registers_reg[27][15]  ( .G(n2047), .D(n2106), .Q(
        \registers[27][15] ) );
  DLH_X1 \registers_reg[27][14]  ( .G(n2047), .D(n2109), .Q(
        \registers[27][14] ) );
  DLH_X1 \registers_reg[27][13]  ( .G(n2047), .D(n2112), .Q(
        \registers[27][13] ) );
  DLH_X1 \registers_reg[27][12]  ( .G(n2047), .D(n2115), .Q(
        \registers[27][12] ) );
  DLH_X1 \registers_reg[27][11]  ( .G(n2048), .D(n2118), .Q(
        \registers[27][11] ) );
  DLH_X1 \registers_reg[27][10]  ( .G(n2048), .D(n2121), .Q(
        \registers[27][10] ) );
  DLH_X1 \registers_reg[27][9]  ( .G(n2048), .D(n2124), .Q(\registers[27][9] )
         );
  DLH_X1 \registers_reg[27][8]  ( .G(n2048), .D(n2127), .Q(\registers[27][8] )
         );
  DLH_X1 \registers_reg[27][7]  ( .G(n2048), .D(n2130), .Q(\registers[27][7] )
         );
  DLH_X1 \registers_reg[27][6]  ( .G(n2048), .D(n2133), .Q(\registers[27][6] )
         );
  DLH_X1 \registers_reg[27][5]  ( .G(n2048), .D(n2136), .Q(\registers[27][5] )
         );
  DLH_X1 \registers_reg[27][4]  ( .G(n2048), .D(n2139), .Q(\registers[27][4] )
         );
  DLH_X1 \registers_reg[27][3]  ( .G(n2048), .D(n2142), .Q(\registers[27][3] )
         );
  DLH_X1 \registers_reg[27][2]  ( .G(n2048), .D(n2145), .Q(\registers[27][2] )
         );
  DLH_X1 \registers_reg[27][1]  ( .G(n2046), .D(n2148), .Q(\registers[27][1] )
         );
  DLH_X1 \registers_reg[27][0]  ( .G(n2046), .D(n2151), .Q(\registers[27][0] )
         );
  DLH_X1 \registers_reg[28][31]  ( .G(n2049), .D(n2058), .Q(
        \registers[28][31] ) );
  DLH_X1 \registers_reg[28][30]  ( .G(n2049), .D(n2061), .Q(
        \registers[28][30] ) );
  DLH_X1 \registers_reg[28][29]  ( .G(n2049), .D(n2064), .Q(
        \registers[28][29] ) );
  DLH_X1 \registers_reg[28][28]  ( .G(n2049), .D(n2067), .Q(
        \registers[28][28] ) );
  DLH_X1 \registers_reg[28][27]  ( .G(n2049), .D(n2070), .Q(
        \registers[28][27] ) );
  DLH_X1 \registers_reg[28][26]  ( .G(n2049), .D(n2073), .Q(
        \registers[28][26] ) );
  DLH_X1 \registers_reg[28][25]  ( .G(n2049), .D(n2076), .Q(
        \registers[28][25] ) );
  DLH_X1 \registers_reg[28][24]  ( .G(n2050), .D(n2079), .Q(
        \registers[28][24] ) );
  DLH_X1 \registers_reg[28][23]  ( .G(n2050), .D(n2082), .Q(
        \registers[28][23] ) );
  DLH_X1 \registers_reg[28][22]  ( .G(n2050), .D(n2085), .Q(
        \registers[28][22] ) );
  DLH_X1 \registers_reg[28][21]  ( .G(n2050), .D(n2088), .Q(
        \registers[28][21] ) );
  DLH_X1 \registers_reg[28][20]  ( .G(n2049), .D(n2091), .Q(
        \registers[28][20] ) );
  DLH_X1 \registers_reg[28][19]  ( .G(n2050), .D(n2094), .Q(
        \registers[28][19] ) );
  DLH_X1 \registers_reg[28][18]  ( .G(n2050), .D(n2097), .Q(
        \registers[28][18] ) );
  DLH_X1 \registers_reg[28][17]  ( .G(n2049), .D(n2100), .Q(
        \registers[28][17] ) );
  DLH_X1 \registers_reg[28][16]  ( .G(n2050), .D(n2103), .Q(
        \registers[28][16] ) );
  DLH_X1 \registers_reg[28][15]  ( .G(n2050), .D(n2106), .Q(
        \registers[28][15] ) );
  DLH_X1 \registers_reg[28][14]  ( .G(n2050), .D(n2109), .Q(
        \registers[28][14] ) );
  DLH_X1 \registers_reg[28][13]  ( .G(n2050), .D(n2112), .Q(
        \registers[28][13] ) );
  DLH_X1 \registers_reg[28][12]  ( .G(n2050), .D(n2115), .Q(
        \registers[28][12] ) );
  DLH_X1 \registers_reg[28][11]  ( .G(n2051), .D(n2118), .Q(
        \registers[28][11] ) );
  DLH_X1 \registers_reg[28][10]  ( .G(n2051), .D(n2121), .Q(
        \registers[28][10] ) );
  DLH_X1 \registers_reg[28][9]  ( .G(n2051), .D(n2124), .Q(\registers[28][9] )
         );
  DLH_X1 \registers_reg[28][8]  ( .G(n2051), .D(n2127), .Q(\registers[28][8] )
         );
  DLH_X1 \registers_reg[28][7]  ( .G(n2051), .D(n2130), .Q(\registers[28][7] )
         );
  DLH_X1 \registers_reg[28][6]  ( .G(n2051), .D(n2133), .Q(\registers[28][6] )
         );
  DLH_X1 \registers_reg[28][5]  ( .G(n2051), .D(n2136), .Q(\registers[28][5] )
         );
  DLH_X1 \registers_reg[28][4]  ( .G(n2051), .D(n2139), .Q(\registers[28][4] )
         );
  DLH_X1 \registers_reg[28][3]  ( .G(n2051), .D(n2142), .Q(\registers[28][3] )
         );
  DLH_X1 \registers_reg[28][2]  ( .G(n2051), .D(n2145), .Q(\registers[28][2] )
         );
  DLH_X1 \registers_reg[28][1]  ( .G(n2049), .D(n2148), .Q(\registers[28][1] )
         );
  DLH_X1 \registers_reg[28][0]  ( .G(n2049), .D(n2151), .Q(\registers[28][0] )
         );
  DLH_X1 \registers_reg[29][31]  ( .G(n2052), .D(n2058), .Q(
        \registers[29][31] ) );
  DLH_X1 \registers_reg[29][30]  ( .G(n2052), .D(n2061), .Q(
        \registers[29][30] ) );
  DLH_X1 \registers_reg[29][29]  ( .G(n2052), .D(n2064), .Q(
        \registers[29][29] ) );
  DLH_X1 \registers_reg[29][28]  ( .G(n2052), .D(n2067), .Q(
        \registers[29][28] ) );
  DLH_X1 \registers_reg[29][27]  ( .G(n2052), .D(n2070), .Q(
        \registers[29][27] ) );
  DLH_X1 \registers_reg[29][26]  ( .G(n2052), .D(n2073), .Q(
        \registers[29][26] ) );
  DLH_X1 \registers_reg[29][25]  ( .G(n2052), .D(n2076), .Q(
        \registers[29][25] ) );
  DLH_X1 \registers_reg[29][24]  ( .G(n2053), .D(n2079), .Q(
        \registers[29][24] ) );
  DLH_X1 \registers_reg[29][23]  ( .G(n2053), .D(n2082), .Q(
        \registers[29][23] ) );
  DLH_X1 \registers_reg[29][22]  ( .G(n2053), .D(n2085), .Q(
        \registers[29][22] ) );
  DLH_X1 \registers_reg[29][21]  ( .G(n2053), .D(n2088), .Q(
        \registers[29][21] ) );
  DLH_X1 \registers_reg[29][20]  ( .G(n2052), .D(n2091), .Q(
        \registers[29][20] ) );
  DLH_X1 \registers_reg[29][19]  ( .G(n2053), .D(n2094), .Q(
        \registers[29][19] ) );
  DLH_X1 \registers_reg[29][18]  ( .G(n2053), .D(n2097), .Q(
        \registers[29][18] ) );
  DLH_X1 \registers_reg[29][17]  ( .G(n2052), .D(n2100), .Q(
        \registers[29][17] ) );
  DLH_X1 \registers_reg[29][16]  ( .G(n2053), .D(n2103), .Q(
        \registers[29][16] ) );
  DLH_X1 \registers_reg[29][15]  ( .G(n2053), .D(n2106), .Q(
        \registers[29][15] ) );
  DLH_X1 \registers_reg[29][14]  ( .G(n2053), .D(n2109), .Q(
        \registers[29][14] ) );
  DLH_X1 \registers_reg[29][13]  ( .G(n2053), .D(n2112), .Q(
        \registers[29][13] ) );
  DLH_X1 \registers_reg[29][12]  ( .G(n2053), .D(n2115), .Q(
        \registers[29][12] ) );
  DLH_X1 \registers_reg[29][11]  ( .G(n2054), .D(n2118), .Q(
        \registers[29][11] ) );
  DLH_X1 \registers_reg[29][10]  ( .G(n2054), .D(n2121), .Q(
        \registers[29][10] ) );
  DLH_X1 \registers_reg[29][9]  ( .G(n2054), .D(n2124), .Q(\registers[29][9] )
         );
  DLH_X1 \registers_reg[29][8]  ( .G(n2054), .D(n2127), .Q(\registers[29][8] )
         );
  DLH_X1 \registers_reg[29][7]  ( .G(n2054), .D(n2130), .Q(\registers[29][7] )
         );
  DLH_X1 \registers_reg[29][6]  ( .G(n2054), .D(n2133), .Q(\registers[29][6] )
         );
  DLH_X1 \registers_reg[29][5]  ( .G(n2054), .D(n2136), .Q(\registers[29][5] )
         );
  DLH_X1 \registers_reg[29][4]  ( .G(n2054), .D(n2139), .Q(\registers[29][4] )
         );
  DLH_X1 \registers_reg[29][3]  ( .G(n2054), .D(n2142), .Q(\registers[29][3] )
         );
  DLH_X1 \registers_reg[29][2]  ( .G(n2054), .D(n2145), .Q(\registers[29][2] )
         );
  DLH_X1 \registers_reg[29][1]  ( .G(n2052), .D(n2148), .Q(\registers[29][1] )
         );
  DLH_X1 \registers_reg[29][0]  ( .G(n2052), .D(n2151), .Q(\registers[29][0] )
         );
  DLH_X1 \registers_reg[30][31]  ( .G(n2055), .D(n2058), .Q(
        \registers[30][31] ) );
  DLH_X1 \registers_reg[30][30]  ( .G(n2055), .D(n2061), .Q(
        \registers[30][30] ) );
  DLH_X1 \registers_reg[30][29]  ( .G(n2055), .D(n2064), .Q(
        \registers[30][29] ) );
  DLH_X1 \registers_reg[30][28]  ( .G(n2055), .D(n2067), .Q(
        \registers[30][28] ) );
  DLH_X1 \registers_reg[30][27]  ( .G(n2055), .D(n2070), .Q(
        \registers[30][27] ) );
  DLH_X1 \registers_reg[30][26]  ( .G(n2055), .D(n2073), .Q(
        \registers[30][26] ) );
  DLH_X1 \registers_reg[30][25]  ( .G(n2055), .D(n2076), .Q(
        \registers[30][25] ) );
  DLH_X1 \registers_reg[30][24]  ( .G(n2056), .D(n2079), .Q(
        \registers[30][24] ) );
  DLH_X1 \registers_reg[30][23]  ( .G(n2056), .D(n2082), .Q(
        \registers[30][23] ) );
  DLH_X1 \registers_reg[30][22]  ( .G(n2056), .D(n2085), .Q(
        \registers[30][22] ) );
  DLH_X1 \registers_reg[30][21]  ( .G(n2056), .D(n2088), .Q(
        \registers[30][21] ) );
  DLH_X1 \registers_reg[30][20]  ( .G(n2055), .D(n2091), .Q(
        \registers[30][20] ) );
  DLH_X1 \registers_reg[30][19]  ( .G(n2056), .D(n2094), .Q(
        \registers[30][19] ) );
  DLH_X1 \registers_reg[30][18]  ( .G(n2056), .D(n2097), .Q(
        \registers[30][18] ) );
  DLH_X1 \registers_reg[30][17]  ( .G(n2055), .D(n2100), .Q(
        \registers[30][17] ) );
  DLH_X1 \registers_reg[30][16]  ( .G(n2056), .D(n2103), .Q(
        \registers[30][16] ) );
  DLH_X1 \registers_reg[30][15]  ( .G(n2056), .D(n2106), .Q(
        \registers[30][15] ) );
  DLH_X1 \registers_reg[30][14]  ( .G(n2056), .D(n2109), .Q(
        \registers[30][14] ) );
  DLH_X1 \registers_reg[30][13]  ( .G(n2056), .D(n2112), .Q(
        \registers[30][13] ) );
  DLH_X1 \registers_reg[30][12]  ( .G(n2056), .D(n2115), .Q(
        \registers[30][12] ) );
  DLH_X1 \registers_reg[30][11]  ( .G(n2057), .D(n2118), .Q(
        \registers[30][11] ) );
  DLH_X1 \registers_reg[30][10]  ( .G(n2057), .D(n2121), .Q(
        \registers[30][10] ) );
  DLH_X1 \registers_reg[30][9]  ( .G(n2057), .D(n2124), .Q(\registers[30][9] )
         );
  DLH_X1 \registers_reg[30][8]  ( .G(n2057), .D(n2127), .Q(\registers[30][8] )
         );
  DLH_X1 \registers_reg[30][7]  ( .G(n2057), .D(n2130), .Q(\registers[30][7] )
         );
  DLH_X1 \registers_reg[30][6]  ( .G(n2057), .D(n2133), .Q(\registers[30][6] )
         );
  DLH_X1 \registers_reg[30][5]  ( .G(n2057), .D(n2136), .Q(\registers[30][5] )
         );
  DLH_X1 \registers_reg[30][4]  ( .G(n2057), .D(n2139), .Q(\registers[30][4] )
         );
  DLH_X1 \registers_reg[30][3]  ( .G(n2057), .D(n2142), .Q(\registers[30][3] )
         );
  DLH_X1 \registers_reg[30][2]  ( .G(n2057), .D(n2145), .Q(\registers[30][2] )
         );
  DLH_X1 \registers_reg[30][1]  ( .G(n2055), .D(n2148), .Q(\registers[30][1] )
         );
  DLH_X1 \registers_reg[30][0]  ( .G(n2055), .D(n2151), .Q(\registers[30][0] )
         );
  DLH_X1 \registers_reg[31][31]  ( .G(n2154), .D(n2058), .Q(
        \registers[31][31] ) );
  DLH_X1 \registers_reg[31][30]  ( .G(n2154), .D(n2061), .Q(
        \registers[31][30] ) );
  DLH_X1 \registers_reg[31][29]  ( .G(n2154), .D(n2064), .Q(
        \registers[31][29] ) );
  DLH_X1 \registers_reg[31][28]  ( .G(n2154), .D(n2067), .Q(
        \registers[31][28] ) );
  DLH_X1 \registers_reg[31][27]  ( .G(n2154), .D(n2070), .Q(
        \registers[31][27] ) );
  DLH_X1 \registers_reg[31][26]  ( .G(n2154), .D(n2073), .Q(
        \registers[31][26] ) );
  DLH_X1 \registers_reg[31][25]  ( .G(n2154), .D(n2076), .Q(
        \registers[31][25] ) );
  DLH_X1 \registers_reg[31][24]  ( .G(n2155), .D(n2079), .Q(
        \registers[31][24] ) );
  DLH_X1 \registers_reg[31][23]  ( .G(n2155), .D(n2082), .Q(
        \registers[31][23] ) );
  DLH_X1 \registers_reg[31][22]  ( .G(n2155), .D(n2085), .Q(
        \registers[31][22] ) );
  DLH_X1 \registers_reg[31][21]  ( .G(n2155), .D(n2088), .Q(
        \registers[31][21] ) );
  DLH_X1 \registers_reg[31][20]  ( .G(n2154), .D(n2091), .Q(
        \registers[31][20] ) );
  DLH_X1 \registers_reg[31][19]  ( .G(n2155), .D(n2094), .Q(
        \registers[31][19] ) );
  DLH_X1 \registers_reg[31][18]  ( .G(n2155), .D(n2097), .Q(
        \registers[31][18] ) );
  DLH_X1 \registers_reg[31][17]  ( .G(n2154), .D(n2100), .Q(
        \registers[31][17] ) );
  DLH_X1 \registers_reg[31][16]  ( .G(n2155), .D(n2103), .Q(
        \registers[31][16] ) );
  DLH_X1 \registers_reg[31][15]  ( .G(n2155), .D(n2106), .Q(
        \registers[31][15] ) );
  DLH_X1 \registers_reg[31][14]  ( .G(n2155), .D(n2109), .Q(
        \registers[31][14] ) );
  DLH_X1 \registers_reg[31][13]  ( .G(n2155), .D(n2112), .Q(
        \registers[31][13] ) );
  DLH_X1 \registers_reg[31][12]  ( .G(n2155), .D(n2115), .Q(
        \registers[31][12] ) );
  DLH_X1 \registers_reg[31][11]  ( .G(n2156), .D(n2118), .Q(
        \registers[31][11] ) );
  DLH_X1 \registers_reg[31][10]  ( .G(n2156), .D(n2121), .Q(
        \registers[31][10] ) );
  DLH_X1 \registers_reg[31][9]  ( .G(n2156), .D(n2124), .Q(\registers[31][9] )
         );
  DLH_X1 \registers_reg[31][8]  ( .G(n2156), .D(n2127), .Q(\registers[31][8] )
         );
  DLH_X1 \registers_reg[31][7]  ( .G(n2156), .D(n2130), .Q(\registers[31][7] )
         );
  DLH_X1 \registers_reg[31][6]  ( .G(n2156), .D(n2133), .Q(\registers[31][6] )
         );
  DLH_X1 \registers_reg[31][5]  ( .G(n2156), .D(n2136), .Q(\registers[31][5] )
         );
  DLH_X1 \registers_reg[31][4]  ( .G(n2156), .D(n2139), .Q(\registers[31][4] )
         );
  DLH_X1 \registers_reg[31][3]  ( .G(n2156), .D(n2142), .Q(\registers[31][3] )
         );
  DLH_X1 \registers_reg[31][2]  ( .G(n2156), .D(n2145), .Q(\registers[31][2] )
         );
  DLH_X1 \registers_reg[31][1]  ( .G(n2154), .D(n2148), .Q(\registers[31][1] )
         );
  DLH_X1 \registers_reg[31][0]  ( .G(n2154), .D(n2151), .Q(\registers[31][0] )
         );
  DLH_X1 \out2_reg[31]  ( .G(n1962), .D(N243), .Q(out2[31]) );
  DLH_X1 \out2_reg[30]  ( .G(n1962), .D(N244), .Q(out2[30]) );
  DLH_X1 \out2_reg[29]  ( .G(n1962), .D(N245), .Q(out2[29]) );
  DLH_X1 \out2_reg[28]  ( .G(n1963), .D(N246), .Q(out2[28]) );
  DLH_X1 \out2_reg[27]  ( .G(n1962), .D(N247), .Q(out2[27]) );
  DLH_X1 \out2_reg[26]  ( .G(n1963), .D(N248), .Q(out2[26]) );
  DLH_X1 \out2_reg[25]  ( .G(n1963), .D(N249), .Q(out2[25]) );
  DLH_X1 \out2_reg[24]  ( .G(n1964), .D(N250), .Q(out2[24]) );
  DLH_X1 \out2_reg[23]  ( .G(n1964), .D(N251), .Q(out2[23]) );
  DLH_X1 \out2_reg[22]  ( .G(n1964), .D(N252), .Q(out2[22]) );
  DLH_X1 \out2_reg[21]  ( .G(n1965), .D(N253), .Q(out2[21]) );
  DLH_X1 \out2_reg[20]  ( .G(n1963), .D(N254), .Q(out2[20]) );
  DLH_X1 \out2_reg[19]  ( .G(n1964), .D(N255), .Q(out2[19]) );
  DLH_X1 \out2_reg[18]  ( .G(n1964), .D(N256), .Q(out2[18]) );
  DLH_X1 \out2_reg[17]  ( .G(n1962), .D(N257), .Q(out2[17]) );
  DLH_X1 \out2_reg[16]  ( .G(n1964), .D(N258), .Q(out2[16]) );
  DLH_X1 \out2_reg[15]  ( .G(n1965), .D(N259), .Q(out2[15]) );
  DLH_X1 \out2_reg[14]  ( .G(n1965), .D(N260), .Q(out2[14]) );
  DLH_X1 \out2_reg[13]  ( .G(n1965), .D(N261), .Q(out2[13]) );
  DLH_X1 \out2_reg[12]  ( .G(n1965), .D(N262), .Q(out2[12]) );
  DLH_X1 \out2_reg[11]  ( .G(n1966), .D(N263), .Q(out2[11]) );
  DLH_X1 \out2_reg[10]  ( .G(n1966), .D(N264), .Q(out2[10]) );
  DLH_X1 \out2_reg[9]  ( .G(n1966), .D(N265), .Q(out2[9]) );
  DLH_X1 \out2_reg[8]  ( .G(n1966), .D(N266), .Q(out2[8]) );
  DLH_X1 \out2_reg[7]  ( .G(n1966), .D(N267), .Q(out2[7]) );
  DLH_X1 \out2_reg[6]  ( .G(n1967), .D(N268), .Q(out2[6]) );
  DLH_X1 \out2_reg[5]  ( .G(n1967), .D(N269), .Q(out2[5]) );
  DLH_X1 \out2_reg[4]  ( .G(n1967), .D(N270), .Q(out2[4]) );
  DLH_X1 \out2_reg[3]  ( .G(n1966), .D(N271), .Q(out2[3]) );
  DLH_X1 \out2_reg[2]  ( .G(n1967), .D(N272), .Q(out2[2]) );
  DLH_X1 \out2_reg[1]  ( .G(n1963), .D(N273), .Q(out2[1]) );
  DLH_X1 \out2_reg[0]  ( .G(n1962), .D(N274), .Q(out2[0]) );
  DLH_X1 \out1_reg[31]  ( .G(n1962), .D(N146), .Q(out1[31]) );
  DLH_X1 \out1_reg[30]  ( .G(n1962), .D(N147), .Q(out1[30]) );
  DLH_X1 \out1_reg[29]  ( .G(n1962), .D(N148), .Q(out1[29]) );
  DLH_X1 \out1_reg[28]  ( .G(n1963), .D(N149), .Q(out1[28]) );
  DLH_X1 \out1_reg[27]  ( .G(n1963), .D(N150), .Q(out1[27]) );
  DLH_X1 \out1_reg[26]  ( .G(n1963), .D(N151), .Q(out1[26]) );
  DLH_X1 \out1_reg[25]  ( .G(n1963), .D(N152), .Q(out1[25]) );
  DLH_X1 \out1_reg[24]  ( .G(n1964), .D(N153), .Q(out1[24]) );
  DLH_X1 \out1_reg[23]  ( .G(n1964), .D(N154), .Q(out1[23]) );
  DLH_X1 \out1_reg[22]  ( .G(n1964), .D(N155), .Q(out1[22]) );
  DLH_X1 \out1_reg[21]  ( .G(n1965), .D(N156), .Q(out1[21]) );
  DLH_X1 \out1_reg[20]  ( .G(n1963), .D(N157), .Q(out1[20]) );
  DLH_X1 \out1_reg[19]  ( .G(n1964), .D(N158), .Q(out1[19]) );
  DLH_X1 \out1_reg[18]  ( .G(n1965), .D(N159), .Q(out1[18]) );
  DLH_X1 \out1_reg[17]  ( .G(n1962), .D(N160), .Q(out1[17]) );
  DLH_X1 \out1_reg[16]  ( .G(n1964), .D(N161), .Q(out1[16]) );
  DLH_X1 \out1_reg[15]  ( .G(n1965), .D(N162), .Q(out1[15]) );
  DLH_X1 \out1_reg[14]  ( .G(n1965), .D(N163), .Q(out1[14]) );
  DLH_X1 \out1_reg[13]  ( .G(n1965), .D(N164), .Q(out1[13]) );
  DLH_X1 \out1_reg[12]  ( .G(n1965), .D(N165), .Q(out1[12]) );
  DLH_X1 \out1_reg[11]  ( .G(n1966), .D(N166), .Q(out1[11]) );
  DLH_X1 \out1_reg[10]  ( .G(n1966), .D(N167), .Q(out1[10]) );
  DLH_X1 \out1_reg[9]  ( .G(n1966), .D(N168), .Q(out1[9]) );
  DLH_X1 \out1_reg[8]  ( .G(n1966), .D(N169), .Q(out1[8]) );
  DLH_X1 \out1_reg[7]  ( .G(n1967), .D(N170), .Q(out1[7]) );
  DLH_X1 \out1_reg[6]  ( .G(n1967), .D(N171), .Q(out1[6]) );
  DLH_X1 \out1_reg[5]  ( .G(n1967), .D(N172), .Q(out1[5]) );
  DLH_X1 \out1_reg[4]  ( .G(n1967), .D(N173), .Q(out1[4]) );
  DLH_X1 \out1_reg[3]  ( .G(n1966), .D(N174), .Q(out1[3]) );
  DLH_X1 \out1_reg[2]  ( .G(n1967), .D(N175), .Q(out1[2]) );
  DLH_X1 \out1_reg[1]  ( .G(n1963), .D(N176), .Q(out1[1]) );
  DLH_X1 \out1_reg[0]  ( .G(n1962), .D(N177), .Q(out1[0]) );
  NAND3_X1 U1832 ( .A1(n2165), .A2(n2164), .A3(n535), .ZN(n527) );
  NAND3_X1 U1833 ( .A1(n535), .A2(n2164), .A3(add_wr[3]), .ZN(n536) );
  NAND3_X1 U1834 ( .A1(n535), .A2(n2165), .A3(add_wr[4]), .ZN(n538) );
  NAND3_X1 U1835 ( .A1(n2167), .A2(n2166), .A3(n2168), .ZN(n537) );
  NAND3_X1 U1836 ( .A1(n2167), .A2(n2166), .A3(add_wr[0]), .ZN(n528) );
  NAND3_X1 U1837 ( .A1(n2168), .A2(n2166), .A3(add_wr[1]), .ZN(n529) );
  NAND3_X1 U1838 ( .A1(add_wr[0]), .A2(n2166), .A3(add_wr[1]), .ZN(n530) );
  NAND3_X1 U1839 ( .A1(n2168), .A2(n2167), .A3(add_wr[2]), .ZN(n531) );
  NAND3_X1 U1840 ( .A1(add_wr[0]), .A2(n2167), .A3(add_wr[2]), .ZN(n532) );
  NAND3_X1 U1841 ( .A1(add_wr[1]), .A2(n2168), .A3(add_wr[2]), .ZN(n533) );
  NAND3_X1 U1842 ( .A1(add_wr[3]), .A2(n535), .A3(add_wr[4]), .ZN(n539) );
  NAND3_X1 U1843 ( .A1(add_wr[1]), .A2(add_wr[0]), .A3(add_wr[2]), .ZN(n534)
         );
  NOR2_X1 U3 ( .A1(n2683), .A2(add_rd1[2]), .ZN(n1697) );
  NOR2_X1 U4 ( .A1(n2687), .A2(add_rd2[2]), .ZN(n1110) );
  BUF_X1 U5 ( .A(n2157), .Z(n2161) );
  BUF_X1 U6 ( .A(n2157), .Z(n2160) );
  BUF_X1 U7 ( .A(n2157), .Z(n2159) );
  BUF_X1 U8 ( .A(n2158), .Z(n2162) );
  BUF_X1 U9 ( .A(n2158), .Z(n2163) );
  BUF_X1 U10 ( .A(reset), .Z(n2157) );
  BUF_X1 U11 ( .A(reset), .Z(n2158) );
  BUF_X1 U12 ( .A(n579), .Z(n1888) );
  BUF_X1 U13 ( .A(n584), .Z(n1876) );
  BUF_X1 U14 ( .A(n579), .Z(n1887) );
  BUF_X1 U15 ( .A(n584), .Z(n1875) );
  BUF_X1 U16 ( .A(n548), .Z(n1960) );
  BUF_X1 U17 ( .A(n553), .Z(n1948) );
  BUF_X1 U18 ( .A(n548), .Z(n1959) );
  BUF_X1 U19 ( .A(n553), .Z(n1947) );
  BUF_X1 U20 ( .A(n551), .Z(n1954) );
  BUF_X1 U21 ( .A(n556), .Z(n1942) );
  BUF_X1 U22 ( .A(n561), .Z(n1930) );
  BUF_X1 U23 ( .A(n566), .Z(n1918) );
  BUF_X1 U24 ( .A(n576), .Z(n1897) );
  BUF_X1 U25 ( .A(n551), .Z(n1953) );
  BUF_X1 U26 ( .A(n556), .Z(n1941) );
  BUF_X1 U27 ( .A(n561), .Z(n1929) );
  BUF_X1 U28 ( .A(n566), .Z(n1917) );
  BUF_X1 U29 ( .A(n576), .Z(n1896) );
  BUF_X1 U30 ( .A(n558), .Z(n1936) );
  BUF_X1 U31 ( .A(n563), .Z(n1924) );
  BUF_X1 U32 ( .A(n573), .Z(n1903) );
  BUF_X1 U33 ( .A(n558), .Z(n1935) );
  BUF_X1 U34 ( .A(n563), .Z(n1923) );
  BUF_X1 U35 ( .A(n573), .Z(n1902) );
  BUF_X1 U36 ( .A(n568), .Z(n1912) );
  BUF_X1 U37 ( .A(n568), .Z(n1911) );
  BUF_X1 U38 ( .A(n552), .Z(n1951) );
  BUF_X1 U39 ( .A(n557), .Z(n1939) );
  BUF_X1 U40 ( .A(n562), .Z(n1927) );
  BUF_X1 U41 ( .A(n567), .Z(n1915) );
  BUF_X1 U42 ( .A(n577), .Z(n1894) );
  BUF_X1 U43 ( .A(n552), .Z(n1950) );
  BUF_X1 U44 ( .A(n557), .Z(n1938) );
  BUF_X1 U45 ( .A(n562), .Z(n1926) );
  BUF_X1 U46 ( .A(n567), .Z(n1914) );
  BUF_X1 U47 ( .A(n577), .Z(n1893) );
  BUF_X1 U48 ( .A(n1158), .Z(n1816) );
  BUF_X1 U49 ( .A(n1158), .Z(n1815) );
  BUF_X1 U50 ( .A(n1168), .Z(n1792) );
  BUF_X1 U51 ( .A(n1173), .Z(n1780) );
  BUF_X1 U52 ( .A(n1168), .Z(n1791) );
  BUF_X1 U53 ( .A(n1173), .Z(n1779) );
  BUF_X1 U54 ( .A(n1169), .Z(n1789) );
  BUF_X1 U55 ( .A(n1174), .Z(n1777) );
  BUF_X1 U56 ( .A(n1169), .Z(n1788) );
  BUF_X1 U57 ( .A(n1174), .Z(n1776) );
  BUF_X1 U58 ( .A(n1159), .Z(n1813) );
  BUF_X1 U59 ( .A(n1159), .Z(n1812) );
  BUF_X1 U60 ( .A(n1161), .Z(n1807) );
  BUF_X1 U61 ( .A(n1161), .Z(n1806) );
  BUF_X1 U62 ( .A(n1136), .Z(n1864) );
  BUF_X1 U63 ( .A(n1141), .Z(n1852) );
  BUF_X1 U64 ( .A(n1146), .Z(n1840) );
  BUF_X1 U65 ( .A(n1151), .Z(n1828) );
  BUF_X1 U66 ( .A(n1136), .Z(n1863) );
  BUF_X1 U67 ( .A(n1141), .Z(n1851) );
  BUF_X1 U68 ( .A(n1146), .Z(n1839) );
  BUF_X1 U69 ( .A(n1151), .Z(n1827) );
  BUF_X1 U70 ( .A(n1165), .Z(n1798) );
  BUF_X1 U71 ( .A(n1170), .Z(n1786) );
  BUF_X1 U72 ( .A(n1165), .Z(n1797) );
  BUF_X1 U73 ( .A(n1170), .Z(n1785) );
  BUF_X1 U74 ( .A(n1155), .Z(n1819) );
  BUF_X1 U75 ( .A(n1155), .Z(n1818) );
  BUF_X1 U76 ( .A(n572), .Z(n1906) );
  BUF_X1 U77 ( .A(n572), .Z(n1905) );
  BUF_X1 U78 ( .A(n582), .Z(n1882) );
  BUF_X1 U79 ( .A(n587), .Z(n1870) );
  BUF_X1 U80 ( .A(n582), .Z(n1881) );
  BUF_X1 U81 ( .A(n587), .Z(n1869) );
  BUF_X1 U82 ( .A(n1138), .Z(n1861) );
  BUF_X1 U83 ( .A(n1143), .Z(n1849) );
  BUF_X1 U84 ( .A(n1148), .Z(n1837) );
  BUF_X1 U85 ( .A(n1153), .Z(n1825) );
  BUF_X1 U86 ( .A(n1163), .Z(n1804) );
  BUF_X1 U87 ( .A(n1138), .Z(n1860) );
  BUF_X1 U88 ( .A(n1143), .Z(n1848) );
  BUF_X1 U89 ( .A(n1148), .Z(n1836) );
  BUF_X1 U90 ( .A(n1153), .Z(n1824) );
  BUF_X1 U91 ( .A(n1163), .Z(n1803) );
  BUF_X1 U92 ( .A(n1166), .Z(n1795) );
  BUF_X1 U93 ( .A(n1171), .Z(n1783) );
  BUF_X1 U94 ( .A(n1166), .Z(n1794) );
  BUF_X1 U95 ( .A(n1171), .Z(n1782) );
  BUF_X1 U96 ( .A(n579), .Z(n1889) );
  BUF_X1 U97 ( .A(n584), .Z(n1877) );
  BUF_X1 U98 ( .A(n578), .Z(n1891) );
  BUF_X1 U99 ( .A(n583), .Z(n1879) );
  BUF_X1 U100 ( .A(n578), .Z(n1890) );
  BUF_X1 U101 ( .A(n583), .Z(n1878) );
  BUF_X1 U102 ( .A(n581), .Z(n1885) );
  BUF_X1 U103 ( .A(n571), .Z(n1909) );
  BUF_X1 U104 ( .A(n581), .Z(n1884) );
  BUF_X1 U105 ( .A(n571), .Z(n1908) );
  BUF_X1 U106 ( .A(n586), .Z(n1873) );
  BUF_X1 U107 ( .A(n586), .Z(n1872) );
  BUF_X1 U108 ( .A(n1160), .Z(n1810) );
  BUF_X1 U109 ( .A(n1160), .Z(n1809) );
  BUF_X1 U110 ( .A(n1135), .Z(n1867) );
  BUF_X1 U111 ( .A(n1140), .Z(n1855) );
  BUF_X1 U112 ( .A(n1145), .Z(n1843) );
  BUF_X1 U113 ( .A(n1150), .Z(n1831) );
  BUF_X1 U114 ( .A(n1135), .Z(n1866) );
  BUF_X1 U115 ( .A(n1140), .Z(n1854) );
  BUF_X1 U116 ( .A(n1145), .Z(n1842) );
  BUF_X1 U117 ( .A(n1150), .Z(n1830) );
  BUF_X1 U118 ( .A(n548), .Z(n1961) );
  BUF_X1 U119 ( .A(n553), .Z(n1949) );
  BUF_X1 U120 ( .A(n551), .Z(n1955) );
  BUF_X1 U121 ( .A(n556), .Z(n1943) );
  BUF_X1 U122 ( .A(n561), .Z(n1931) );
  BUF_X1 U123 ( .A(n566), .Z(n1919) );
  BUF_X1 U124 ( .A(n576), .Z(n1898) );
  BUF_X1 U125 ( .A(n558), .Z(n1937) );
  BUF_X1 U126 ( .A(n563), .Z(n1925) );
  BUF_X1 U127 ( .A(n573), .Z(n1904) );
  BUF_X1 U128 ( .A(n568), .Z(n1913) );
  BUF_X1 U129 ( .A(n552), .Z(n1952) );
  BUF_X1 U130 ( .A(n557), .Z(n1940) );
  BUF_X1 U131 ( .A(n562), .Z(n1928) );
  BUF_X1 U132 ( .A(n567), .Z(n1916) );
  BUF_X1 U133 ( .A(n577), .Z(n1895) );
  BUF_X1 U134 ( .A(n1158), .Z(n1817) );
  BUF_X1 U135 ( .A(n1168), .Z(n1793) );
  BUF_X1 U136 ( .A(n1173), .Z(n1781) );
  BUF_X1 U137 ( .A(n1169), .Z(n1790) );
  BUF_X1 U138 ( .A(n1174), .Z(n1778) );
  BUF_X1 U139 ( .A(n1159), .Z(n1814) );
  BUF_X1 U140 ( .A(n549), .Z(n1957) );
  BUF_X1 U141 ( .A(n549), .Z(n1956) );
  BUF_X1 U142 ( .A(n554), .Z(n1945) );
  BUF_X1 U143 ( .A(n564), .Z(n1921) );
  BUF_X1 U144 ( .A(n554), .Z(n1944) );
  BUF_X1 U145 ( .A(n564), .Z(n1920) );
  BUF_X1 U146 ( .A(n559), .Z(n1933) );
  BUF_X1 U147 ( .A(n574), .Z(n1900) );
  BUF_X1 U148 ( .A(n559), .Z(n1932) );
  BUF_X1 U149 ( .A(n574), .Z(n1899) );
  BUF_X1 U150 ( .A(n1139), .Z(n1857) );
  BUF_X1 U151 ( .A(n1144), .Z(n1845) );
  BUF_X1 U152 ( .A(n1149), .Z(n1833) );
  BUF_X1 U153 ( .A(n1154), .Z(n1821) );
  BUF_X1 U154 ( .A(n1164), .Z(n1800) );
  BUF_X1 U155 ( .A(n1139), .Z(n1858) );
  BUF_X1 U156 ( .A(n1144), .Z(n1846) );
  BUF_X1 U157 ( .A(n1149), .Z(n1834) );
  BUF_X1 U158 ( .A(n1154), .Z(n1822) );
  BUF_X1 U159 ( .A(n1164), .Z(n1801) );
  BUF_X1 U160 ( .A(n1161), .Z(n1808) );
  BUF_X1 U161 ( .A(n1136), .Z(n1865) );
  BUF_X1 U162 ( .A(n1141), .Z(n1853) );
  BUF_X1 U163 ( .A(n1151), .Z(n1829) );
  BUF_X1 U164 ( .A(n1146), .Z(n1841) );
  BUF_X1 U165 ( .A(n1165), .Z(n1799) );
  BUF_X1 U166 ( .A(n1170), .Z(n1787) );
  BUF_X1 U167 ( .A(n1155), .Z(n1820) );
  BUF_X1 U168 ( .A(n572), .Z(n1907) );
  BUF_X1 U169 ( .A(n582), .Z(n1883) );
  BUF_X1 U170 ( .A(n587), .Z(n1871) );
  BUF_X1 U171 ( .A(n1138), .Z(n1862) );
  BUF_X1 U172 ( .A(n1143), .Z(n1850) );
  BUF_X1 U173 ( .A(n1148), .Z(n1838) );
  BUF_X1 U174 ( .A(n1153), .Z(n1826) );
  BUF_X1 U175 ( .A(n1163), .Z(n1805) );
  BUF_X1 U176 ( .A(n1166), .Z(n1796) );
  BUF_X1 U177 ( .A(n1171), .Z(n1784) );
  BUF_X1 U178 ( .A(n578), .Z(n1892) );
  BUF_X1 U179 ( .A(n583), .Z(n1880) );
  BUF_X1 U180 ( .A(n581), .Z(n1886) );
  BUF_X1 U181 ( .A(n571), .Z(n1910) );
  BUF_X1 U182 ( .A(n586), .Z(n1874) );
  BUF_X1 U183 ( .A(n1160), .Z(n1811) );
  BUF_X1 U184 ( .A(n1135), .Z(n1868) );
  BUF_X1 U185 ( .A(n1140), .Z(n1856) );
  BUF_X1 U186 ( .A(n1145), .Z(n1844) );
  BUF_X1 U187 ( .A(n1150), .Z(n1832) );
  BUF_X1 U188 ( .A(n549), .Z(n1958) );
  BUF_X1 U189 ( .A(n554), .Z(n1946) );
  BUF_X1 U190 ( .A(n564), .Z(n1922) );
  BUF_X1 U191 ( .A(n559), .Z(n1934) );
  BUF_X1 U192 ( .A(n574), .Z(n1901) );
  BUF_X1 U193 ( .A(n1139), .Z(n1859) );
  BUF_X1 U194 ( .A(n1144), .Z(n1847) );
  BUF_X1 U195 ( .A(n1149), .Z(n1835) );
  BUF_X1 U196 ( .A(n1154), .Z(n1823) );
  BUF_X1 U197 ( .A(n1164), .Z(n1802) );
  BUF_X1 U198 ( .A(N307), .Z(n2155) );
  BUF_X1 U199 ( .A(N307), .Z(n2154) );
  BUF_X1 U200 ( .A(N340), .Z(n2056) );
  BUF_X1 U201 ( .A(N340), .Z(n2055) );
  BUF_X1 U202 ( .A(N341), .Z(n2053) );
  BUF_X1 U203 ( .A(N341), .Z(n2052) );
  BUF_X1 U204 ( .A(N342), .Z(n2050) );
  BUF_X1 U205 ( .A(N342), .Z(n2049) );
  BUF_X1 U206 ( .A(N343), .Z(n2047) );
  BUF_X1 U207 ( .A(N343), .Z(n2046) );
  BUF_X1 U208 ( .A(N344), .Z(n2044) );
  BUF_X1 U209 ( .A(N344), .Z(n2043) );
  BUF_X1 U210 ( .A(N345), .Z(n2041) );
  BUF_X1 U211 ( .A(N345), .Z(n2040) );
  BUF_X1 U212 ( .A(N346), .Z(n2038) );
  BUF_X1 U213 ( .A(N346), .Z(n2037) );
  BUF_X1 U214 ( .A(N347), .Z(n2035) );
  BUF_X1 U215 ( .A(N347), .Z(n2034) );
  BUF_X1 U216 ( .A(N348), .Z(n2032) );
  BUF_X1 U217 ( .A(N348), .Z(n2031) );
  BUF_X1 U218 ( .A(N349), .Z(n2029) );
  BUF_X1 U219 ( .A(N349), .Z(n2028) );
  BUF_X1 U220 ( .A(N350), .Z(n2026) );
  BUF_X1 U221 ( .A(N350), .Z(n2025) );
  BUF_X1 U222 ( .A(N351), .Z(n2023) );
  BUF_X1 U223 ( .A(N351), .Z(n2022) );
  BUF_X1 U224 ( .A(N352), .Z(n2020) );
  BUF_X1 U225 ( .A(N352), .Z(n2019) );
  BUF_X1 U226 ( .A(N353), .Z(n2017) );
  BUF_X1 U227 ( .A(N353), .Z(n2016) );
  BUF_X1 U228 ( .A(N354), .Z(n2014) );
  BUF_X1 U229 ( .A(N354), .Z(n2013) );
  BUF_X1 U230 ( .A(N355), .Z(n2011) );
  BUF_X1 U231 ( .A(N355), .Z(n2010) );
  BUF_X1 U232 ( .A(N356), .Z(n2008) );
  BUF_X1 U233 ( .A(N356), .Z(n2007) );
  BUF_X1 U234 ( .A(N357), .Z(n2005) );
  BUF_X1 U235 ( .A(N357), .Z(n2004) );
  BUF_X1 U236 ( .A(N358), .Z(n2002) );
  BUF_X1 U237 ( .A(N358), .Z(n2001) );
  BUF_X1 U238 ( .A(N359), .Z(n1998) );
  BUF_X1 U239 ( .A(N359), .Z(n1999) );
  BUF_X1 U240 ( .A(N360), .Z(n1995) );
  BUF_X1 U241 ( .A(N360), .Z(n1996) );
  BUF_X1 U242 ( .A(N361), .Z(n1992) );
  BUF_X1 U243 ( .A(N361), .Z(n1993) );
  BUF_X1 U244 ( .A(N362), .Z(n1989) );
  BUF_X1 U245 ( .A(N362), .Z(n1990) );
  BUF_X1 U246 ( .A(N363), .Z(n1986) );
  BUF_X1 U247 ( .A(N363), .Z(n1987) );
  BUF_X1 U248 ( .A(N364), .Z(n1983) );
  BUF_X1 U249 ( .A(N364), .Z(n1984) );
  BUF_X1 U250 ( .A(N365), .Z(n1980) );
  BUF_X1 U251 ( .A(N365), .Z(n1981) );
  BUF_X1 U252 ( .A(N366), .Z(n1977) );
  BUF_X1 U253 ( .A(N366), .Z(n1978) );
  BUF_X1 U254 ( .A(N367), .Z(n1974) );
  BUF_X1 U255 ( .A(N367), .Z(n1975) );
  BUF_X1 U256 ( .A(N368), .Z(n1971) );
  BUF_X1 U257 ( .A(N368), .Z(n1972) );
  BUF_X1 U258 ( .A(N369), .Z(n1968) );
  BUF_X1 U259 ( .A(N369), .Z(n1969) );
  BUF_X1 U260 ( .A(N308), .Z(n2151) );
  BUF_X1 U261 ( .A(N316), .Z(n2127) );
  BUF_X1 U262 ( .A(N317), .Z(n2124) );
  BUF_X1 U263 ( .A(N318), .Z(n2121) );
  BUF_X1 U264 ( .A(N319), .Z(n2118) );
  BUF_X1 U265 ( .A(N320), .Z(n2115) );
  BUF_X1 U266 ( .A(N321), .Z(n2112) );
  BUF_X1 U267 ( .A(N322), .Z(n2109) );
  BUF_X1 U268 ( .A(N323), .Z(n2106) );
  BUF_X1 U269 ( .A(N324), .Z(n2103) );
  BUF_X1 U270 ( .A(N325), .Z(n2100) );
  BUF_X1 U271 ( .A(N326), .Z(n2097) );
  BUF_X1 U272 ( .A(N327), .Z(n2094) );
  BUF_X1 U273 ( .A(N328), .Z(n2091) );
  BUF_X1 U274 ( .A(N329), .Z(n2088) );
  BUF_X1 U275 ( .A(N330), .Z(n2085) );
  BUF_X1 U276 ( .A(N331), .Z(n2082) );
  BUF_X1 U277 ( .A(N332), .Z(n2079) );
  BUF_X1 U278 ( .A(N333), .Z(n2076) );
  BUF_X1 U279 ( .A(N334), .Z(n2073) );
  BUF_X1 U280 ( .A(N335), .Z(n2070) );
  BUF_X1 U281 ( .A(N336), .Z(n2067) );
  BUF_X1 U282 ( .A(N337), .Z(n2064) );
  BUF_X1 U283 ( .A(N338), .Z(n2061) );
  BUF_X1 U284 ( .A(N339), .Z(n2058) );
  BUF_X1 U285 ( .A(N308), .Z(n2152) );
  BUF_X1 U286 ( .A(N316), .Z(n2128) );
  BUF_X1 U287 ( .A(N317), .Z(n2125) );
  BUF_X1 U288 ( .A(N318), .Z(n2122) );
  BUF_X1 U289 ( .A(N319), .Z(n2119) );
  BUF_X1 U290 ( .A(N320), .Z(n2116) );
  BUF_X1 U291 ( .A(N321), .Z(n2113) );
  BUF_X1 U292 ( .A(N322), .Z(n2110) );
  BUF_X1 U293 ( .A(N323), .Z(n2107) );
  BUF_X1 U294 ( .A(N324), .Z(n2104) );
  BUF_X1 U295 ( .A(N325), .Z(n2101) );
  BUF_X1 U296 ( .A(N326), .Z(n2098) );
  BUF_X1 U297 ( .A(N327), .Z(n2095) );
  BUF_X1 U298 ( .A(N328), .Z(n2092) );
  BUF_X1 U299 ( .A(N329), .Z(n2089) );
  BUF_X1 U300 ( .A(N330), .Z(n2086) );
  BUF_X1 U301 ( .A(N331), .Z(n2083) );
  BUF_X1 U302 ( .A(N332), .Z(n2080) );
  BUF_X1 U303 ( .A(N333), .Z(n2077) );
  BUF_X1 U304 ( .A(N334), .Z(n2074) );
  BUF_X1 U305 ( .A(N335), .Z(n2071) );
  BUF_X1 U306 ( .A(N336), .Z(n2068) );
  BUF_X1 U307 ( .A(N337), .Z(n2065) );
  BUF_X1 U308 ( .A(N338), .Z(n2062) );
  BUF_X1 U309 ( .A(N339), .Z(n2059) );
  BUF_X1 U310 ( .A(N309), .Z(n2148) );
  BUF_X1 U311 ( .A(N310), .Z(n2145) );
  BUF_X1 U312 ( .A(N311), .Z(n2142) );
  BUF_X1 U313 ( .A(N312), .Z(n2139) );
  BUF_X1 U314 ( .A(N313), .Z(n2136) );
  BUF_X1 U315 ( .A(N314), .Z(n2133) );
  BUF_X1 U316 ( .A(N315), .Z(n2130) );
  BUF_X1 U317 ( .A(N309), .Z(n2149) );
  BUF_X1 U318 ( .A(N310), .Z(n2146) );
  BUF_X1 U319 ( .A(N311), .Z(n2143) );
  BUF_X1 U320 ( .A(N312), .Z(n2140) );
  BUF_X1 U321 ( .A(N313), .Z(n2137) );
  BUF_X1 U322 ( .A(N314), .Z(n2134) );
  BUF_X1 U323 ( .A(N315), .Z(n2131) );
  BUF_X1 U324 ( .A(N307), .Z(n2156) );
  BUF_X1 U325 ( .A(N340), .Z(n2057) );
  BUF_X1 U326 ( .A(N341), .Z(n2054) );
  BUF_X1 U327 ( .A(N342), .Z(n2051) );
  BUF_X1 U328 ( .A(N343), .Z(n2048) );
  BUF_X1 U329 ( .A(N344), .Z(n2045) );
  BUF_X1 U330 ( .A(N345), .Z(n2042) );
  BUF_X1 U331 ( .A(N346), .Z(n2039) );
  BUF_X1 U332 ( .A(N347), .Z(n2036) );
  BUF_X1 U333 ( .A(N348), .Z(n2033) );
  BUF_X1 U334 ( .A(N349), .Z(n2030) );
  BUF_X1 U335 ( .A(N350), .Z(n2027) );
  BUF_X1 U336 ( .A(N351), .Z(n2024) );
  BUF_X1 U337 ( .A(N352), .Z(n2021) );
  BUF_X1 U338 ( .A(N353), .Z(n2018) );
  BUF_X1 U339 ( .A(N354), .Z(n2015) );
  BUF_X1 U340 ( .A(N355), .Z(n2012) );
  BUF_X1 U341 ( .A(N356), .Z(n2009) );
  BUF_X1 U342 ( .A(N357), .Z(n2006) );
  BUF_X1 U343 ( .A(N358), .Z(n2003) );
  BUF_X1 U344 ( .A(N359), .Z(n2000) );
  BUF_X1 U345 ( .A(N360), .Z(n1997) );
  BUF_X1 U346 ( .A(N361), .Z(n1994) );
  BUF_X1 U347 ( .A(N362), .Z(n1991) );
  BUF_X1 U348 ( .A(N363), .Z(n1988) );
  BUF_X1 U349 ( .A(N364), .Z(n1985) );
  BUF_X1 U350 ( .A(N365), .Z(n1982) );
  BUF_X1 U351 ( .A(N366), .Z(n1979) );
  BUF_X1 U352 ( .A(N367), .Z(n1976) );
  BUF_X1 U353 ( .A(N368), .Z(n1973) );
  BUF_X1 U354 ( .A(N369), .Z(n1970) );
  BUF_X1 U355 ( .A(N308), .Z(n2153) );
  BUF_X1 U356 ( .A(N316), .Z(n2129) );
  BUF_X1 U357 ( .A(N317), .Z(n2126) );
  BUF_X1 U358 ( .A(N318), .Z(n2123) );
  BUF_X1 U359 ( .A(N319), .Z(n2120) );
  BUF_X1 U360 ( .A(N320), .Z(n2117) );
  BUF_X1 U361 ( .A(N321), .Z(n2114) );
  BUF_X1 U362 ( .A(N322), .Z(n2111) );
  BUF_X1 U363 ( .A(N323), .Z(n2108) );
  BUF_X1 U364 ( .A(N324), .Z(n2105) );
  BUF_X1 U365 ( .A(N325), .Z(n2102) );
  BUF_X1 U366 ( .A(N326), .Z(n2099) );
  BUF_X1 U367 ( .A(N327), .Z(n2096) );
  BUF_X1 U368 ( .A(N328), .Z(n2093) );
  BUF_X1 U369 ( .A(N329), .Z(n2090) );
  BUF_X1 U370 ( .A(N330), .Z(n2087) );
  BUF_X1 U371 ( .A(N331), .Z(n2084) );
  BUF_X1 U372 ( .A(N332), .Z(n2081) );
  BUF_X1 U373 ( .A(N333), .Z(n2078) );
  BUF_X1 U374 ( .A(N334), .Z(n2075) );
  BUF_X1 U375 ( .A(N335), .Z(n2072) );
  BUF_X1 U376 ( .A(N336), .Z(n2069) );
  BUF_X1 U377 ( .A(N337), .Z(n2066) );
  BUF_X1 U378 ( .A(N338), .Z(n2063) );
  BUF_X1 U379 ( .A(N339), .Z(n2060) );
  BUF_X1 U380 ( .A(N309), .Z(n2150) );
  BUF_X1 U381 ( .A(N310), .Z(n2147) );
  BUF_X1 U382 ( .A(N311), .Z(n2144) );
  BUF_X1 U383 ( .A(N312), .Z(n2141) );
  BUF_X1 U384 ( .A(N313), .Z(n2138) );
  BUF_X1 U385 ( .A(N314), .Z(n2135) );
  BUF_X1 U386 ( .A(N315), .Z(n2132) );
  NOR2_X1 U387 ( .A1(n2683), .A2(n2682), .ZN(n1699) );
  NOR2_X1 U388 ( .A1(n2687), .A2(n2686), .ZN(n1112) );
  NOR4_X1 U389 ( .A1(n1298), .A2(n1299), .A3(n1300), .A4(n1301), .ZN(n1297) );
  OAI221_X1 U390 ( .B1(n2672), .B2(n1831), .C1(n2640), .C2(n1828), .A(n1305), 
        .ZN(n1298) );
  OAI221_X1 U391 ( .B1(n2608), .B2(n1843), .C1(n2576), .C2(n1840), .A(n1304), 
        .ZN(n1299) );
  OAI221_X1 U392 ( .B1(n2544), .B2(n1855), .C1(n2512), .C2(n1852), .A(n1303), 
        .ZN(n1300) );
  NOR4_X1 U393 ( .A1(n1315), .A2(n1316), .A3(n1317), .A4(n1318), .ZN(n1314) );
  OAI221_X1 U394 ( .B1(n2671), .B2(n1831), .C1(n2639), .C2(n1828), .A(n1322), 
        .ZN(n1315) );
  OAI221_X1 U395 ( .B1(n2607), .B2(n1843), .C1(n2575), .C2(n1840), .A(n1321), 
        .ZN(n1316) );
  OAI221_X1 U396 ( .B1(n2543), .B2(n1855), .C1(n2511), .C2(n1852), .A(n1320), 
        .ZN(n1317) );
  NOR4_X1 U397 ( .A1(n1332), .A2(n1333), .A3(n1334), .A4(n1335), .ZN(n1331) );
  OAI221_X1 U398 ( .B1(n2670), .B2(n1831), .C1(n2638), .C2(n1828), .A(n1339), 
        .ZN(n1332) );
  OAI221_X1 U399 ( .B1(n2606), .B2(n1843), .C1(n2574), .C2(n1840), .A(n1338), 
        .ZN(n1333) );
  OAI221_X1 U400 ( .B1(n2542), .B2(n1855), .C1(n2510), .C2(n1852), .A(n1337), 
        .ZN(n1334) );
  NOR4_X1 U401 ( .A1(n1349), .A2(n1350), .A3(n1351), .A4(n1352), .ZN(n1348) );
  OAI221_X1 U402 ( .B1(n2669), .B2(n1831), .C1(n2637), .C2(n1828), .A(n1356), 
        .ZN(n1349) );
  OAI221_X1 U403 ( .B1(n2605), .B2(n1843), .C1(n2573), .C2(n1840), .A(n1355), 
        .ZN(n1350) );
  OAI221_X1 U404 ( .B1(n2541), .B2(n1855), .C1(n2509), .C2(n1852), .A(n1354), 
        .ZN(n1351) );
  NOR4_X1 U405 ( .A1(n1366), .A2(n1367), .A3(n1368), .A4(n1369), .ZN(n1365) );
  OAI221_X1 U406 ( .B1(n2668), .B2(n1831), .C1(n2636), .C2(n1828), .A(n1373), 
        .ZN(n1366) );
  OAI221_X1 U407 ( .B1(n2604), .B2(n1843), .C1(n2572), .C2(n1840), .A(n1372), 
        .ZN(n1367) );
  OAI221_X1 U408 ( .B1(n2540), .B2(n1855), .C1(n2508), .C2(n1852), .A(n1371), 
        .ZN(n1368) );
  NOR4_X1 U409 ( .A1(n1383), .A2(n1384), .A3(n1385), .A4(n1386), .ZN(n1382) );
  OAI221_X1 U410 ( .B1(n2667), .B2(n1831), .C1(n2635), .C2(n1828), .A(n1390), 
        .ZN(n1383) );
  OAI221_X1 U411 ( .B1(n2603), .B2(n1843), .C1(n2571), .C2(n1840), .A(n1389), 
        .ZN(n1384) );
  OAI221_X1 U412 ( .B1(n2539), .B2(n1855), .C1(n2507), .C2(n1852), .A(n1388), 
        .ZN(n1385) );
  NOR4_X1 U413 ( .A1(n1400), .A2(n1401), .A3(n1402), .A4(n1403), .ZN(n1399) );
  OAI221_X1 U414 ( .B1(n2666), .B2(n1831), .C1(n2634), .C2(n1828), .A(n1407), 
        .ZN(n1400) );
  OAI221_X1 U415 ( .B1(n2602), .B2(n1843), .C1(n2570), .C2(n1840), .A(n1406), 
        .ZN(n1401) );
  OAI221_X1 U416 ( .B1(n2538), .B2(n1855), .C1(n2506), .C2(n1852), .A(n1405), 
        .ZN(n1402) );
  NOR4_X1 U417 ( .A1(n1417), .A2(n1418), .A3(n1419), .A4(n1420), .ZN(n1416) );
  OAI221_X1 U418 ( .B1(n2665), .B2(n1831), .C1(n2633), .C2(n1828), .A(n1424), 
        .ZN(n1417) );
  OAI221_X1 U419 ( .B1(n2601), .B2(n1843), .C1(n2569), .C2(n1840), .A(n1423), 
        .ZN(n1418) );
  OAI221_X1 U420 ( .B1(n2537), .B2(n1855), .C1(n2505), .C2(n1852), .A(n1422), 
        .ZN(n1419) );
  NOR4_X1 U421 ( .A1(n1434), .A2(n1435), .A3(n1436), .A4(n1437), .ZN(n1433) );
  OAI221_X1 U422 ( .B1(n2664), .B2(n1831), .C1(n2632), .C2(n1828), .A(n1441), 
        .ZN(n1434) );
  OAI221_X1 U423 ( .B1(n2600), .B2(n1843), .C1(n2568), .C2(n1840), .A(n1440), 
        .ZN(n1435) );
  OAI221_X1 U424 ( .B1(n2536), .B2(n1855), .C1(n2504), .C2(n1852), .A(n1439), 
        .ZN(n1436) );
  NOR4_X1 U425 ( .A1(n1451), .A2(n1452), .A3(n1453), .A4(n1454), .ZN(n1450) );
  OAI221_X1 U426 ( .B1(n2663), .B2(n1831), .C1(n2631), .C2(n1828), .A(n1458), 
        .ZN(n1451) );
  OAI221_X1 U427 ( .B1(n2599), .B2(n1843), .C1(n2567), .C2(n1840), .A(n1457), 
        .ZN(n1452) );
  OAI221_X1 U428 ( .B1(n2535), .B2(n1855), .C1(n2503), .C2(n1852), .A(n1456), 
        .ZN(n1453) );
  NOR4_X1 U429 ( .A1(n1468), .A2(n1469), .A3(n1470), .A4(n1471), .ZN(n1467) );
  OAI221_X1 U430 ( .B1(n2662), .B2(n1831), .C1(n2630), .C2(n1828), .A(n1475), 
        .ZN(n1468) );
  OAI221_X1 U431 ( .B1(n2598), .B2(n1843), .C1(n2566), .C2(n1840), .A(n1474), 
        .ZN(n1469) );
  OAI221_X1 U432 ( .B1(n2534), .B2(n1855), .C1(n2502), .C2(n1852), .A(n1473), 
        .ZN(n1470) );
  NOR4_X1 U433 ( .A1(n1485), .A2(n1486), .A3(n1487), .A4(n1488), .ZN(n1484) );
  OAI221_X1 U434 ( .B1(n2661), .B2(n1831), .C1(n2629), .C2(n1828), .A(n1492), 
        .ZN(n1485) );
  OAI221_X1 U435 ( .B1(n2597), .B2(n1843), .C1(n2565), .C2(n1840), .A(n1491), 
        .ZN(n1486) );
  OAI221_X1 U436 ( .B1(n2533), .B2(n1855), .C1(n2501), .C2(n1852), .A(n1490), 
        .ZN(n1487) );
  NOR4_X1 U437 ( .A1(n1502), .A2(n1503), .A3(n1504), .A4(n1505), .ZN(n1501) );
  OAI221_X1 U438 ( .B1(n2660), .B2(n1830), .C1(n2628), .C2(n1827), .A(n1509), 
        .ZN(n1502) );
  OAI221_X1 U439 ( .B1(n2596), .B2(n1842), .C1(n2564), .C2(n1839), .A(n1508), 
        .ZN(n1503) );
  OAI221_X1 U440 ( .B1(n2532), .B2(n1854), .C1(n2500), .C2(n1851), .A(n1507), 
        .ZN(n1504) );
  NOR4_X1 U441 ( .A1(n1519), .A2(n1520), .A3(n1521), .A4(n1522), .ZN(n1518) );
  OAI221_X1 U442 ( .B1(n2659), .B2(n1830), .C1(n2627), .C2(n1827), .A(n1526), 
        .ZN(n1519) );
  OAI221_X1 U443 ( .B1(n2595), .B2(n1842), .C1(n2563), .C2(n1839), .A(n1525), 
        .ZN(n1520) );
  OAI221_X1 U444 ( .B1(n2531), .B2(n1854), .C1(n2499), .C2(n1851), .A(n1524), 
        .ZN(n1521) );
  NOR4_X1 U445 ( .A1(n1536), .A2(n1537), .A3(n1538), .A4(n1539), .ZN(n1535) );
  OAI221_X1 U446 ( .B1(n2658), .B2(n1830), .C1(n2626), .C2(n1827), .A(n1543), 
        .ZN(n1536) );
  OAI221_X1 U447 ( .B1(n2594), .B2(n1842), .C1(n2562), .C2(n1839), .A(n1542), 
        .ZN(n1537) );
  OAI221_X1 U448 ( .B1(n2530), .B2(n1854), .C1(n2498), .C2(n1851), .A(n1541), 
        .ZN(n1538) );
  NOR4_X1 U449 ( .A1(n1553), .A2(n1554), .A3(n1555), .A4(n1556), .ZN(n1552) );
  OAI221_X1 U450 ( .B1(n2657), .B2(n1830), .C1(n2625), .C2(n1827), .A(n1560), 
        .ZN(n1553) );
  OAI221_X1 U451 ( .B1(n2593), .B2(n1842), .C1(n2561), .C2(n1839), .A(n1559), 
        .ZN(n1554) );
  OAI221_X1 U452 ( .B1(n2529), .B2(n1854), .C1(n2497), .C2(n1851), .A(n1558), 
        .ZN(n1555) );
  NOR4_X1 U453 ( .A1(n1570), .A2(n1571), .A3(n1572), .A4(n1573), .ZN(n1569) );
  OAI221_X1 U454 ( .B1(n2656), .B2(n1830), .C1(n2624), .C2(n1827), .A(n1577), 
        .ZN(n1570) );
  OAI221_X1 U455 ( .B1(n2592), .B2(n1842), .C1(n2560), .C2(n1839), .A(n1576), 
        .ZN(n1571) );
  OAI221_X1 U456 ( .B1(n2528), .B2(n1854), .C1(n2496), .C2(n1851), .A(n1575), 
        .ZN(n1572) );
  NOR4_X1 U457 ( .A1(n1587), .A2(n1588), .A3(n1589), .A4(n1590), .ZN(n1586) );
  OAI221_X1 U458 ( .B1(n2655), .B2(n1830), .C1(n2623), .C2(n1827), .A(n1594), 
        .ZN(n1587) );
  OAI221_X1 U459 ( .B1(n2591), .B2(n1842), .C1(n2559), .C2(n1839), .A(n1593), 
        .ZN(n1588) );
  OAI221_X1 U460 ( .B1(n2527), .B2(n1854), .C1(n2495), .C2(n1851), .A(n1592), 
        .ZN(n1589) );
  NOR4_X1 U461 ( .A1(n1604), .A2(n1605), .A3(n1606), .A4(n1607), .ZN(n1603) );
  OAI221_X1 U462 ( .B1(n2654), .B2(n1830), .C1(n2622), .C2(n1827), .A(n1611), 
        .ZN(n1604) );
  OAI221_X1 U463 ( .B1(n2590), .B2(n1842), .C1(n2558), .C2(n1839), .A(n1610), 
        .ZN(n1605) );
  OAI221_X1 U464 ( .B1(n2526), .B2(n1854), .C1(n2494), .C2(n1851), .A(n1609), 
        .ZN(n1606) );
  NOR4_X1 U465 ( .A1(n1621), .A2(n1622), .A3(n1623), .A4(n1624), .ZN(n1620) );
  OAI221_X1 U466 ( .B1(n2653), .B2(n1830), .C1(n2621), .C2(n1827), .A(n1628), 
        .ZN(n1621) );
  OAI221_X1 U467 ( .B1(n2589), .B2(n1842), .C1(n2557), .C2(n1839), .A(n1627), 
        .ZN(n1622) );
  OAI221_X1 U468 ( .B1(n2525), .B2(n1854), .C1(n2493), .C2(n1851), .A(n1626), 
        .ZN(n1623) );
  NOR4_X1 U469 ( .A1(n1638), .A2(n1639), .A3(n1640), .A4(n1641), .ZN(n1637) );
  OAI221_X1 U470 ( .B1(n2652), .B2(n1830), .C1(n2620), .C2(n1827), .A(n1645), 
        .ZN(n1638) );
  OAI221_X1 U471 ( .B1(n2588), .B2(n1842), .C1(n2556), .C2(n1839), .A(n1644), 
        .ZN(n1639) );
  OAI221_X1 U472 ( .B1(n2524), .B2(n1854), .C1(n2492), .C2(n1851), .A(n1643), 
        .ZN(n1640) );
  NOR4_X1 U473 ( .A1(n1655), .A2(n1656), .A3(n1657), .A4(n1658), .ZN(n1654) );
  OAI221_X1 U474 ( .B1(n2651), .B2(n1830), .C1(n2619), .C2(n1827), .A(n1662), 
        .ZN(n1655) );
  OAI221_X1 U475 ( .B1(n2587), .B2(n1842), .C1(n2555), .C2(n1839), .A(n1661), 
        .ZN(n1656) );
  OAI221_X1 U476 ( .B1(n2523), .B2(n1854), .C1(n2491), .C2(n1851), .A(n1660), 
        .ZN(n1657) );
  NOR4_X1 U477 ( .A1(n1672), .A2(n1673), .A3(n1674), .A4(n1675), .ZN(n1671) );
  OAI221_X1 U478 ( .B1(n2650), .B2(n1830), .C1(n2618), .C2(n1827), .A(n1679), 
        .ZN(n1672) );
  OAI221_X1 U479 ( .B1(n2586), .B2(n1842), .C1(n2554), .C2(n1839), .A(n1678), 
        .ZN(n1673) );
  OAI221_X1 U480 ( .B1(n2522), .B2(n1854), .C1(n2490), .C2(n1851), .A(n1677), 
        .ZN(n1674) );
  NOR4_X1 U481 ( .A1(n1689), .A2(n1690), .A3(n1691), .A4(n1692), .ZN(n1688) );
  OAI221_X1 U482 ( .B1(n2649), .B2(n1830), .C1(n2617), .C2(n1827), .A(n1704), 
        .ZN(n1689) );
  OAI221_X1 U483 ( .B1(n2585), .B2(n1842), .C1(n2553), .C2(n1839), .A(n1701), 
        .ZN(n1690) );
  OAI221_X1 U484 ( .B1(n2521), .B2(n1854), .C1(n2489), .C2(n1851), .A(n1698), 
        .ZN(n1691) );
  NOR4_X1 U485 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1130) );
  OAI221_X1 U486 ( .B1(n2680), .B2(n1832), .C1(n2648), .C2(n1829), .A(n1152), 
        .ZN(n1131) );
  OAI221_X1 U487 ( .B1(n2616), .B2(n1844), .C1(n2584), .C2(n1841), .A(n1147), 
        .ZN(n1132) );
  OAI221_X1 U488 ( .B1(n2552), .B2(n1856), .C1(n2520), .C2(n1853), .A(n1142), 
        .ZN(n1133) );
  NOR4_X1 U489 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1178) );
  OAI221_X1 U490 ( .B1(n2679), .B2(n1832), .C1(n2647), .C2(n1829), .A(n1186), 
        .ZN(n1179) );
  OAI221_X1 U491 ( .B1(n2615), .B2(n1844), .C1(n2583), .C2(n1841), .A(n1185), 
        .ZN(n1180) );
  OAI221_X1 U492 ( .B1(n2551), .B2(n1856), .C1(n2519), .C2(n1853), .A(n1184), 
        .ZN(n1181) );
  NOR4_X1 U493 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1195) );
  OAI221_X1 U494 ( .B1(n2678), .B2(n1832), .C1(n2646), .C2(n1829), .A(n1203), 
        .ZN(n1196) );
  OAI221_X1 U495 ( .B1(n2614), .B2(n1844), .C1(n2582), .C2(n1841), .A(n1202), 
        .ZN(n1197) );
  OAI221_X1 U496 ( .B1(n2550), .B2(n1856), .C1(n2518), .C2(n1853), .A(n1201), 
        .ZN(n1198) );
  NOR4_X1 U497 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1212) );
  OAI221_X1 U498 ( .B1(n2677), .B2(n1832), .C1(n2645), .C2(n1829), .A(n1220), 
        .ZN(n1213) );
  OAI221_X1 U499 ( .B1(n2613), .B2(n1844), .C1(n2581), .C2(n1841), .A(n1219), 
        .ZN(n1214) );
  OAI221_X1 U500 ( .B1(n2549), .B2(n1856), .C1(n2517), .C2(n1853), .A(n1218), 
        .ZN(n1215) );
  NOR4_X1 U501 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1229) );
  OAI221_X1 U502 ( .B1(n2676), .B2(n1832), .C1(n2644), .C2(n1829), .A(n1237), 
        .ZN(n1230) );
  OAI221_X1 U503 ( .B1(n2612), .B2(n1844), .C1(n2580), .C2(n1841), .A(n1236), 
        .ZN(n1231) );
  OAI221_X1 U504 ( .B1(n2548), .B2(n1856), .C1(n2516), .C2(n1853), .A(n1235), 
        .ZN(n1232) );
  NOR4_X1 U505 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246) );
  OAI221_X1 U506 ( .B1(n2675), .B2(n1832), .C1(n2643), .C2(n1829), .A(n1254), 
        .ZN(n1247) );
  OAI221_X1 U507 ( .B1(n2611), .B2(n1844), .C1(n2579), .C2(n1841), .A(n1253), 
        .ZN(n1248) );
  OAI221_X1 U508 ( .B1(n2547), .B2(n1856), .C1(n2515), .C2(n1853), .A(n1252), 
        .ZN(n1249) );
  NOR4_X1 U509 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1263) );
  OAI221_X1 U510 ( .B1(n2674), .B2(n1832), .C1(n2642), .C2(n1829), .A(n1271), 
        .ZN(n1264) );
  OAI221_X1 U511 ( .B1(n2610), .B2(n1844), .C1(n2578), .C2(n1841), .A(n1270), 
        .ZN(n1265) );
  OAI221_X1 U512 ( .B1(n2546), .B2(n1856), .C1(n2514), .C2(n1853), .A(n1269), 
        .ZN(n1266) );
  NOR4_X1 U513 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1280) );
  OAI221_X1 U514 ( .B1(n2673), .B2(n1832), .C1(n2641), .C2(n1829), .A(n1288), 
        .ZN(n1281) );
  OAI221_X1 U515 ( .B1(n2609), .B2(n1844), .C1(n2577), .C2(n1841), .A(n1287), 
        .ZN(n1282) );
  OAI221_X1 U516 ( .B1(n2545), .B2(n1856), .C1(n2513), .C2(n1853), .A(n1286), 
        .ZN(n1283) );
  NOR4_X1 U517 ( .A1(n544), .A2(n545), .A3(n546), .A4(n547), .ZN(n543) );
  OAI221_X1 U518 ( .B1(n1925), .B2(n2680), .C1(n1922), .C2(n2648), .A(n565), 
        .ZN(n544) );
  OAI221_X1 U519 ( .B1(n1937), .B2(n2616), .C1(n1934), .C2(n2584), .A(n560), 
        .ZN(n545) );
  OAI221_X1 U520 ( .B1(n1949), .B2(n2552), .C1(n1946), .C2(n2520), .A(n555), 
        .ZN(n546) );
  NOR4_X1 U521 ( .A1(n592), .A2(n593), .A3(n594), .A4(n595), .ZN(n591) );
  OAI221_X1 U522 ( .B1(n1925), .B2(n2679), .C1(n1922), .C2(n2647), .A(n599), 
        .ZN(n592) );
  OAI221_X1 U523 ( .B1(n1937), .B2(n2615), .C1(n1934), .C2(n2583), .A(n598), 
        .ZN(n593) );
  OAI221_X1 U524 ( .B1(n1949), .B2(n2551), .C1(n1946), .C2(n2519), .A(n597), 
        .ZN(n594) );
  NOR4_X1 U525 ( .A1(n609), .A2(n610), .A3(n611), .A4(n612), .ZN(n608) );
  OAI221_X1 U526 ( .B1(n1925), .B2(n2678), .C1(n1922), .C2(n2646), .A(n616), 
        .ZN(n609) );
  OAI221_X1 U527 ( .B1(n1937), .B2(n2614), .C1(n1934), .C2(n2582), .A(n615), 
        .ZN(n610) );
  OAI221_X1 U528 ( .B1(n1949), .B2(n2550), .C1(n1946), .C2(n2518), .A(n614), 
        .ZN(n611) );
  NOR4_X1 U529 ( .A1(n626), .A2(n627), .A3(n628), .A4(n629), .ZN(n625) );
  OAI221_X1 U530 ( .B1(n1925), .B2(n2677), .C1(n1922), .C2(n2645), .A(n633), 
        .ZN(n626) );
  OAI221_X1 U531 ( .B1(n1937), .B2(n2613), .C1(n1934), .C2(n2581), .A(n632), 
        .ZN(n627) );
  OAI221_X1 U532 ( .B1(n1949), .B2(n2549), .C1(n1946), .C2(n2517), .A(n631), 
        .ZN(n628) );
  NOR4_X1 U533 ( .A1(n643), .A2(n644), .A3(n645), .A4(n646), .ZN(n642) );
  OAI221_X1 U534 ( .B1(n1925), .B2(n2676), .C1(n1922), .C2(n2644), .A(n650), 
        .ZN(n643) );
  OAI221_X1 U535 ( .B1(n1937), .B2(n2612), .C1(n1934), .C2(n2580), .A(n649), 
        .ZN(n644) );
  OAI221_X1 U536 ( .B1(n1949), .B2(n2548), .C1(n1946), .C2(n2516), .A(n648), 
        .ZN(n645) );
  NOR4_X1 U537 ( .A1(n660), .A2(n661), .A3(n662), .A4(n663), .ZN(n659) );
  OAI221_X1 U538 ( .B1(n1925), .B2(n2675), .C1(n1922), .C2(n2643), .A(n667), 
        .ZN(n660) );
  OAI221_X1 U539 ( .B1(n1937), .B2(n2611), .C1(n1934), .C2(n2579), .A(n666), 
        .ZN(n661) );
  OAI221_X1 U540 ( .B1(n1949), .B2(n2547), .C1(n1946), .C2(n2515), .A(n665), 
        .ZN(n662) );
  NOR4_X1 U541 ( .A1(n677), .A2(n678), .A3(n679), .A4(n680), .ZN(n676) );
  OAI221_X1 U542 ( .B1(n1925), .B2(n2674), .C1(n1922), .C2(n2642), .A(n684), 
        .ZN(n677) );
  OAI221_X1 U543 ( .B1(n1937), .B2(n2610), .C1(n1934), .C2(n2578), .A(n683), 
        .ZN(n678) );
  OAI221_X1 U544 ( .B1(n1949), .B2(n2546), .C1(n1946), .C2(n2514), .A(n682), 
        .ZN(n679) );
  NOR4_X1 U545 ( .A1(n694), .A2(n695), .A3(n696), .A4(n697), .ZN(n693) );
  OAI221_X1 U546 ( .B1(n1925), .B2(n2673), .C1(n1922), .C2(n2641), .A(n701), 
        .ZN(n694) );
  OAI221_X1 U547 ( .B1(n1937), .B2(n2609), .C1(n1934), .C2(n2577), .A(n700), 
        .ZN(n695) );
  OAI221_X1 U548 ( .B1(n1949), .B2(n2545), .C1(n1946), .C2(n2513), .A(n699), 
        .ZN(n696) );
  NOR4_X1 U549 ( .A1(n711), .A2(n712), .A3(n713), .A4(n714), .ZN(n710) );
  OAI221_X1 U550 ( .B1(n1924), .B2(n2672), .C1(n1921), .C2(n2640), .A(n718), 
        .ZN(n711) );
  OAI221_X1 U551 ( .B1(n1936), .B2(n2608), .C1(n1933), .C2(n2576), .A(n717), 
        .ZN(n712) );
  OAI221_X1 U552 ( .B1(n1948), .B2(n2544), .C1(n1945), .C2(n2512), .A(n716), 
        .ZN(n713) );
  NOR4_X1 U553 ( .A1(n728), .A2(n729), .A3(n730), .A4(n731), .ZN(n727) );
  OAI221_X1 U554 ( .B1(n1924), .B2(n2671), .C1(n1921), .C2(n2639), .A(n735), 
        .ZN(n728) );
  OAI221_X1 U555 ( .B1(n1936), .B2(n2607), .C1(n1933), .C2(n2575), .A(n734), 
        .ZN(n729) );
  OAI221_X1 U556 ( .B1(n1948), .B2(n2543), .C1(n1945), .C2(n2511), .A(n733), 
        .ZN(n730) );
  NOR4_X1 U557 ( .A1(n745), .A2(n746), .A3(n747), .A4(n748), .ZN(n744) );
  OAI221_X1 U558 ( .B1(n1924), .B2(n2670), .C1(n1921), .C2(n2638), .A(n752), 
        .ZN(n745) );
  OAI221_X1 U559 ( .B1(n1936), .B2(n2606), .C1(n1933), .C2(n2574), .A(n751), 
        .ZN(n746) );
  OAI221_X1 U560 ( .B1(n1948), .B2(n2542), .C1(n1945), .C2(n2510), .A(n750), 
        .ZN(n747) );
  NOR4_X1 U561 ( .A1(n762), .A2(n763), .A3(n764), .A4(n765), .ZN(n761) );
  OAI221_X1 U562 ( .B1(n1924), .B2(n2669), .C1(n1921), .C2(n2637), .A(n769), 
        .ZN(n762) );
  OAI221_X1 U563 ( .B1(n1936), .B2(n2605), .C1(n1933), .C2(n2573), .A(n768), 
        .ZN(n763) );
  OAI221_X1 U564 ( .B1(n1948), .B2(n2541), .C1(n1945), .C2(n2509), .A(n767), 
        .ZN(n764) );
  NOR4_X1 U565 ( .A1(n779), .A2(n780), .A3(n781), .A4(n782), .ZN(n778) );
  OAI221_X1 U566 ( .B1(n1924), .B2(n2668), .C1(n1921), .C2(n2636), .A(n786), 
        .ZN(n779) );
  OAI221_X1 U567 ( .B1(n1936), .B2(n2604), .C1(n1933), .C2(n2572), .A(n785), 
        .ZN(n780) );
  OAI221_X1 U568 ( .B1(n1948), .B2(n2540), .C1(n1945), .C2(n2508), .A(n784), 
        .ZN(n781) );
  NOR4_X1 U569 ( .A1(n796), .A2(n797), .A3(n798), .A4(n799), .ZN(n795) );
  OAI221_X1 U570 ( .B1(n1924), .B2(n2667), .C1(n1921), .C2(n2635), .A(n803), 
        .ZN(n796) );
  OAI221_X1 U571 ( .B1(n1936), .B2(n2603), .C1(n1933), .C2(n2571), .A(n802), 
        .ZN(n797) );
  OAI221_X1 U572 ( .B1(n1948), .B2(n2539), .C1(n1945), .C2(n2507), .A(n801), 
        .ZN(n798) );
  NOR4_X1 U573 ( .A1(n813), .A2(n814), .A3(n815), .A4(n816), .ZN(n812) );
  OAI221_X1 U574 ( .B1(n1924), .B2(n2666), .C1(n1921), .C2(n2634), .A(n820), 
        .ZN(n813) );
  OAI221_X1 U575 ( .B1(n1936), .B2(n2602), .C1(n1933), .C2(n2570), .A(n819), 
        .ZN(n814) );
  OAI221_X1 U576 ( .B1(n1948), .B2(n2538), .C1(n1945), .C2(n2506), .A(n818), 
        .ZN(n815) );
  NOR4_X1 U577 ( .A1(n830), .A2(n831), .A3(n832), .A4(n833), .ZN(n829) );
  OAI221_X1 U578 ( .B1(n1924), .B2(n2665), .C1(n1921), .C2(n2633), .A(n837), 
        .ZN(n830) );
  OAI221_X1 U579 ( .B1(n1936), .B2(n2601), .C1(n1933), .C2(n2569), .A(n836), 
        .ZN(n831) );
  OAI221_X1 U580 ( .B1(n1948), .B2(n2537), .C1(n1945), .C2(n2505), .A(n835), 
        .ZN(n832) );
  NOR4_X1 U581 ( .A1(n847), .A2(n848), .A3(n849), .A4(n850), .ZN(n846) );
  OAI221_X1 U582 ( .B1(n1924), .B2(n2664), .C1(n1921), .C2(n2632), .A(n854), 
        .ZN(n847) );
  OAI221_X1 U583 ( .B1(n1936), .B2(n2600), .C1(n1933), .C2(n2568), .A(n853), 
        .ZN(n848) );
  OAI221_X1 U584 ( .B1(n1948), .B2(n2536), .C1(n1945), .C2(n2504), .A(n852), 
        .ZN(n849) );
  NOR4_X1 U585 ( .A1(n864), .A2(n865), .A3(n866), .A4(n867), .ZN(n863) );
  OAI221_X1 U586 ( .B1(n1924), .B2(n2663), .C1(n1921), .C2(n2631), .A(n871), 
        .ZN(n864) );
  OAI221_X1 U587 ( .B1(n1936), .B2(n2599), .C1(n1933), .C2(n2567), .A(n870), 
        .ZN(n865) );
  OAI221_X1 U588 ( .B1(n1948), .B2(n2535), .C1(n1945), .C2(n2503), .A(n869), 
        .ZN(n866) );
  NOR4_X1 U589 ( .A1(n881), .A2(n882), .A3(n883), .A4(n884), .ZN(n880) );
  OAI221_X1 U590 ( .B1(n1924), .B2(n2662), .C1(n1921), .C2(n2630), .A(n888), 
        .ZN(n881) );
  OAI221_X1 U591 ( .B1(n1936), .B2(n2598), .C1(n1933), .C2(n2566), .A(n887), 
        .ZN(n882) );
  OAI221_X1 U592 ( .B1(n1948), .B2(n2534), .C1(n1945), .C2(n2502), .A(n886), 
        .ZN(n883) );
  NOR4_X1 U593 ( .A1(n898), .A2(n899), .A3(n900), .A4(n901), .ZN(n897) );
  OAI221_X1 U594 ( .B1(n1924), .B2(n2661), .C1(n1921), .C2(n2629), .A(n905), 
        .ZN(n898) );
  OAI221_X1 U595 ( .B1(n1936), .B2(n2597), .C1(n1933), .C2(n2565), .A(n904), 
        .ZN(n899) );
  OAI221_X1 U596 ( .B1(n1948), .B2(n2533), .C1(n1945), .C2(n2501), .A(n903), 
        .ZN(n900) );
  NOR4_X1 U597 ( .A1(n915), .A2(n916), .A3(n917), .A4(n918), .ZN(n914) );
  OAI221_X1 U598 ( .B1(n1923), .B2(n2660), .C1(n1920), .C2(n2628), .A(n922), 
        .ZN(n915) );
  OAI221_X1 U599 ( .B1(n1935), .B2(n2596), .C1(n1932), .C2(n2564), .A(n921), 
        .ZN(n916) );
  OAI221_X1 U600 ( .B1(n1947), .B2(n2532), .C1(n1944), .C2(n2500), .A(n920), 
        .ZN(n917) );
  NOR4_X1 U601 ( .A1(n932), .A2(n933), .A3(n934), .A4(n935), .ZN(n931) );
  OAI221_X1 U602 ( .B1(n1923), .B2(n2659), .C1(n1920), .C2(n2627), .A(n939), 
        .ZN(n932) );
  OAI221_X1 U603 ( .B1(n1935), .B2(n2595), .C1(n1932), .C2(n2563), .A(n938), 
        .ZN(n933) );
  OAI221_X1 U604 ( .B1(n1947), .B2(n2531), .C1(n1944), .C2(n2499), .A(n937), 
        .ZN(n934) );
  NOR4_X1 U605 ( .A1(n949), .A2(n950), .A3(n951), .A4(n952), .ZN(n948) );
  OAI221_X1 U606 ( .B1(n1923), .B2(n2658), .C1(n1920), .C2(n2626), .A(n956), 
        .ZN(n949) );
  OAI221_X1 U607 ( .B1(n1935), .B2(n2594), .C1(n1932), .C2(n2562), .A(n955), 
        .ZN(n950) );
  OAI221_X1 U608 ( .B1(n1947), .B2(n2530), .C1(n1944), .C2(n2498), .A(n954), 
        .ZN(n951) );
  NOR4_X1 U609 ( .A1(n966), .A2(n967), .A3(n968), .A4(n969), .ZN(n965) );
  OAI221_X1 U610 ( .B1(n1923), .B2(n2657), .C1(n1920), .C2(n2625), .A(n973), 
        .ZN(n966) );
  OAI221_X1 U611 ( .B1(n1935), .B2(n2593), .C1(n1932), .C2(n2561), .A(n972), 
        .ZN(n967) );
  OAI221_X1 U612 ( .B1(n1947), .B2(n2529), .C1(n1944), .C2(n2497), .A(n971), 
        .ZN(n968) );
  NOR4_X1 U613 ( .A1(n983), .A2(n984), .A3(n985), .A4(n986), .ZN(n982) );
  OAI221_X1 U614 ( .B1(n1923), .B2(n2656), .C1(n1920), .C2(n2624), .A(n990), 
        .ZN(n983) );
  OAI221_X1 U615 ( .B1(n1935), .B2(n2592), .C1(n1932), .C2(n2560), .A(n989), 
        .ZN(n984) );
  OAI221_X1 U616 ( .B1(n1947), .B2(n2528), .C1(n1944), .C2(n2496), .A(n988), 
        .ZN(n985) );
  NOR4_X1 U617 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n999) );
  OAI221_X1 U618 ( .B1(n1923), .B2(n2655), .C1(n1920), .C2(n2623), .A(n1007), 
        .ZN(n1000) );
  OAI221_X1 U619 ( .B1(n1935), .B2(n2591), .C1(n1932), .C2(n2559), .A(n1006), 
        .ZN(n1001) );
  OAI221_X1 U620 ( .B1(n1947), .B2(n2527), .C1(n1944), .C2(n2495), .A(n1005), 
        .ZN(n1002) );
  NOR4_X1 U621 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
  OAI221_X1 U622 ( .B1(n1923), .B2(n2654), .C1(n1920), .C2(n2622), .A(n1024), 
        .ZN(n1017) );
  OAI221_X1 U623 ( .B1(n1935), .B2(n2590), .C1(n1932), .C2(n2558), .A(n1023), 
        .ZN(n1018) );
  OAI221_X1 U624 ( .B1(n1947), .B2(n2526), .C1(n1944), .C2(n2494), .A(n1022), 
        .ZN(n1019) );
  NOR4_X1 U625 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1033) );
  OAI221_X1 U626 ( .B1(n1923), .B2(n2653), .C1(n1920), .C2(n2621), .A(n1041), 
        .ZN(n1034) );
  OAI221_X1 U627 ( .B1(n1935), .B2(n2589), .C1(n1932), .C2(n2557), .A(n1040), 
        .ZN(n1035) );
  OAI221_X1 U628 ( .B1(n1947), .B2(n2525), .C1(n1944), .C2(n2493), .A(n1039), 
        .ZN(n1036) );
  NOR4_X1 U629 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
  OAI221_X1 U630 ( .B1(n1923), .B2(n2652), .C1(n1920), .C2(n2620), .A(n1058), 
        .ZN(n1051) );
  OAI221_X1 U631 ( .B1(n1935), .B2(n2588), .C1(n1932), .C2(n2556), .A(n1057), 
        .ZN(n1052) );
  OAI221_X1 U632 ( .B1(n1947), .B2(n2524), .C1(n1944), .C2(n2492), .A(n1056), 
        .ZN(n1053) );
  NOR4_X1 U633 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
  OAI221_X1 U634 ( .B1(n1923), .B2(n2651), .C1(n1920), .C2(n2619), .A(n1075), 
        .ZN(n1068) );
  OAI221_X1 U635 ( .B1(n1935), .B2(n2587), .C1(n1932), .C2(n2555), .A(n1074), 
        .ZN(n1069) );
  OAI221_X1 U636 ( .B1(n1947), .B2(n2523), .C1(n1944), .C2(n2491), .A(n1073), 
        .ZN(n1070) );
  NOR4_X1 U637 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
  OAI221_X1 U638 ( .B1(n1923), .B2(n2650), .C1(n1920), .C2(n2618), .A(n1092), 
        .ZN(n1085) );
  OAI221_X1 U639 ( .B1(n1935), .B2(n2586), .C1(n1932), .C2(n2554), .A(n1091), 
        .ZN(n1086) );
  OAI221_X1 U640 ( .B1(n1947), .B2(n2522), .C1(n1944), .C2(n2490), .A(n1090), 
        .ZN(n1087) );
  NOR4_X1 U641 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1101) );
  OAI221_X1 U642 ( .B1(n1923), .B2(n2649), .C1(n1920), .C2(n2617), .A(n1117), 
        .ZN(n1102) );
  OAI221_X1 U643 ( .B1(n1935), .B2(n2585), .C1(n1932), .C2(n2553), .A(n1114), 
        .ZN(n1103) );
  OAI221_X1 U644 ( .B1(n1947), .B2(n2521), .C1(n1944), .C2(n2489), .A(n1111), 
        .ZN(n1104) );
  OAI22_X1 U645 ( .A1(n1886), .A2(n2392), .B1(n1883), .B2(n2296), .ZN(n580) );
  OAI22_X1 U646 ( .A1(n1874), .A2(n2328), .B1(n1871), .B2(n2424), .ZN(n585) );
  OAI22_X1 U647 ( .A1(n1886), .A2(n2391), .B1(n1883), .B2(n2295), .ZN(n603) );
  OAI22_X1 U648 ( .A1(n1874), .A2(n2327), .B1(n1871), .B2(n2423), .ZN(n604) );
  OAI22_X1 U649 ( .A1(n1886), .A2(n2390), .B1(n1883), .B2(n2294), .ZN(n620) );
  OAI22_X1 U650 ( .A1(n1874), .A2(n2326), .B1(n1871), .B2(n2422), .ZN(n621) );
  OAI22_X1 U651 ( .A1(n1886), .A2(n2389), .B1(n1883), .B2(n2293), .ZN(n637) );
  OAI22_X1 U652 ( .A1(n1874), .A2(n2325), .B1(n1871), .B2(n2421), .ZN(n638) );
  OAI22_X1 U653 ( .A1(n1886), .A2(n2388), .B1(n1883), .B2(n2292), .ZN(n654) );
  OAI22_X1 U654 ( .A1(n1874), .A2(n2324), .B1(n1871), .B2(n2420), .ZN(n655) );
  OAI22_X1 U655 ( .A1(n1886), .A2(n2387), .B1(n1883), .B2(n2291), .ZN(n671) );
  OAI22_X1 U656 ( .A1(n1874), .A2(n2323), .B1(n1871), .B2(n2419), .ZN(n672) );
  OAI22_X1 U657 ( .A1(n1886), .A2(n2386), .B1(n1883), .B2(n2290), .ZN(n688) );
  OAI22_X1 U658 ( .A1(n1874), .A2(n2322), .B1(n1871), .B2(n2418), .ZN(n689) );
  OAI22_X1 U659 ( .A1(n1886), .A2(n2385), .B1(n1883), .B2(n2289), .ZN(n705) );
  OAI22_X1 U660 ( .A1(n1874), .A2(n2321), .B1(n1871), .B2(n2417), .ZN(n706) );
  OAI22_X1 U661 ( .A1(n1910), .A2(n2360), .B1(n1907), .B2(n2232), .ZN(n570) );
  OAI22_X1 U662 ( .A1(n1910), .A2(n2359), .B1(n1907), .B2(n2231), .ZN(n601) );
  OAI22_X1 U663 ( .A1(n1910), .A2(n2358), .B1(n1907), .B2(n2230), .ZN(n618) );
  OAI22_X1 U664 ( .A1(n1910), .A2(n2357), .B1(n1907), .B2(n2229), .ZN(n635) );
  OAI22_X1 U665 ( .A1(n1910), .A2(n2356), .B1(n1907), .B2(n2228), .ZN(n652) );
  OAI22_X1 U666 ( .A1(n1910), .A2(n2355), .B1(n1907), .B2(n2227), .ZN(n669) );
  OAI22_X1 U667 ( .A1(n1910), .A2(n2354), .B1(n1907), .B2(n2226), .ZN(n686) );
  OAI22_X1 U668 ( .A1(n1910), .A2(n2353), .B1(n1907), .B2(n2225), .ZN(n703) );
  OAI22_X1 U669 ( .A1(n2392), .A2(n1793), .B1(n2296), .B2(n1790), .ZN(n1167)
         );
  OAI22_X1 U670 ( .A1(n2328), .A2(n1781), .B1(n2424), .B2(n1778), .ZN(n1172)
         );
  OAI22_X1 U671 ( .A1(n2391), .A2(n1793), .B1(n2295), .B2(n1790), .ZN(n1190)
         );
  OAI22_X1 U672 ( .A1(n2327), .A2(n1781), .B1(n2423), .B2(n1778), .ZN(n1191)
         );
  OAI22_X1 U673 ( .A1(n2390), .A2(n1793), .B1(n2294), .B2(n1790), .ZN(n1207)
         );
  OAI22_X1 U674 ( .A1(n2326), .A2(n1781), .B1(n2422), .B2(n1778), .ZN(n1208)
         );
  OAI22_X1 U675 ( .A1(n2389), .A2(n1793), .B1(n2293), .B2(n1790), .ZN(n1224)
         );
  OAI22_X1 U676 ( .A1(n2325), .A2(n1781), .B1(n2421), .B2(n1778), .ZN(n1225)
         );
  OAI22_X1 U677 ( .A1(n2388), .A2(n1793), .B1(n2292), .B2(n1790), .ZN(n1241)
         );
  OAI22_X1 U678 ( .A1(n2324), .A2(n1781), .B1(n2420), .B2(n1778), .ZN(n1242)
         );
  OAI22_X1 U679 ( .A1(n2387), .A2(n1793), .B1(n2291), .B2(n1790), .ZN(n1258)
         );
  OAI22_X1 U680 ( .A1(n2323), .A2(n1781), .B1(n2419), .B2(n1778), .ZN(n1259)
         );
  OAI22_X1 U681 ( .A1(n2386), .A2(n1793), .B1(n2290), .B2(n1790), .ZN(n1275)
         );
  OAI22_X1 U682 ( .A1(n2322), .A2(n1781), .B1(n2418), .B2(n1778), .ZN(n1276)
         );
  OAI22_X1 U683 ( .A1(n2385), .A2(n1793), .B1(n2289), .B2(n1790), .ZN(n1292)
         );
  OAI22_X1 U684 ( .A1(n2321), .A2(n1781), .B1(n2417), .B2(n1778), .ZN(n1293)
         );
  OAI22_X1 U685 ( .A1(n2360), .A2(n1817), .B1(n2232), .B2(n1814), .ZN(n1157)
         );
  OAI22_X1 U686 ( .A1(n2359), .A2(n1817), .B1(n2231), .B2(n1814), .ZN(n1188)
         );
  OAI22_X1 U687 ( .A1(n2358), .A2(n1817), .B1(n2230), .B2(n1814), .ZN(n1205)
         );
  OAI22_X1 U688 ( .A1(n2357), .A2(n1817), .B1(n2229), .B2(n1814), .ZN(n1222)
         );
  OAI22_X1 U689 ( .A1(n2356), .A2(n1817), .B1(n2228), .B2(n1814), .ZN(n1239)
         );
  OAI22_X1 U690 ( .A1(n2355), .A2(n1817), .B1(n2227), .B2(n1814), .ZN(n1256)
         );
  OAI22_X1 U691 ( .A1(n2354), .A2(n1817), .B1(n2226), .B2(n1814), .ZN(n1273)
         );
  OAI22_X1 U692 ( .A1(n2353), .A2(n1817), .B1(n2225), .B2(n1814), .ZN(n1290)
         );
  OAI22_X1 U693 ( .A1(n2384), .A2(n1792), .B1(n2288), .B2(n1789), .ZN(n1309)
         );
  OAI22_X1 U694 ( .A1(n2320), .A2(n1780), .B1(n2416), .B2(n1777), .ZN(n1310)
         );
  OAI22_X1 U695 ( .A1(n2383), .A2(n1792), .B1(n2287), .B2(n1789), .ZN(n1326)
         );
  OAI22_X1 U696 ( .A1(n2319), .A2(n1780), .B1(n2415), .B2(n1777), .ZN(n1327)
         );
  OAI22_X1 U697 ( .A1(n2382), .A2(n1792), .B1(n2286), .B2(n1789), .ZN(n1343)
         );
  OAI22_X1 U698 ( .A1(n2318), .A2(n1780), .B1(n2414), .B2(n1777), .ZN(n1344)
         );
  OAI22_X1 U699 ( .A1(n2381), .A2(n1792), .B1(n2285), .B2(n1789), .ZN(n1360)
         );
  OAI22_X1 U700 ( .A1(n2317), .A2(n1780), .B1(n2413), .B2(n1777), .ZN(n1361)
         );
  OAI22_X1 U701 ( .A1(n2380), .A2(n1792), .B1(n2284), .B2(n1789), .ZN(n1377)
         );
  OAI22_X1 U702 ( .A1(n2316), .A2(n1780), .B1(n2412), .B2(n1777), .ZN(n1378)
         );
  OAI22_X1 U703 ( .A1(n2379), .A2(n1792), .B1(n2283), .B2(n1789), .ZN(n1394)
         );
  OAI22_X1 U704 ( .A1(n2315), .A2(n1780), .B1(n2411), .B2(n1777), .ZN(n1395)
         );
  OAI22_X1 U705 ( .A1(n2378), .A2(n1792), .B1(n2282), .B2(n1789), .ZN(n1411)
         );
  OAI22_X1 U706 ( .A1(n2314), .A2(n1780), .B1(n2410), .B2(n1777), .ZN(n1412)
         );
  OAI22_X1 U707 ( .A1(n2377), .A2(n1792), .B1(n2281), .B2(n1789), .ZN(n1428)
         );
  OAI22_X1 U708 ( .A1(n2313), .A2(n1780), .B1(n2409), .B2(n1777), .ZN(n1429)
         );
  OAI22_X1 U709 ( .A1(n2376), .A2(n1792), .B1(n2280), .B2(n1789), .ZN(n1445)
         );
  OAI22_X1 U710 ( .A1(n2312), .A2(n1780), .B1(n2408), .B2(n1777), .ZN(n1446)
         );
  OAI22_X1 U711 ( .A1(n2375), .A2(n1792), .B1(n2279), .B2(n1789), .ZN(n1462)
         );
  OAI22_X1 U712 ( .A1(n2311), .A2(n1780), .B1(n2407), .B2(n1777), .ZN(n1463)
         );
  OAI22_X1 U713 ( .A1(n2374), .A2(n1792), .B1(n2278), .B2(n1789), .ZN(n1479)
         );
  OAI22_X1 U714 ( .A1(n2310), .A2(n1780), .B1(n2406), .B2(n1777), .ZN(n1480)
         );
  OAI22_X1 U715 ( .A1(n2373), .A2(n1792), .B1(n2277), .B2(n1789), .ZN(n1496)
         );
  OAI22_X1 U716 ( .A1(n2309), .A2(n1780), .B1(n2405), .B2(n1777), .ZN(n1497)
         );
  OAI22_X1 U717 ( .A1(n2372), .A2(n1791), .B1(n2276), .B2(n1788), .ZN(n1513)
         );
  OAI22_X1 U718 ( .A1(n2308), .A2(n1779), .B1(n2404), .B2(n1776), .ZN(n1514)
         );
  OAI22_X1 U719 ( .A1(n2371), .A2(n1791), .B1(n2275), .B2(n1788), .ZN(n1530)
         );
  OAI22_X1 U720 ( .A1(n2307), .A2(n1779), .B1(n2403), .B2(n1776), .ZN(n1531)
         );
  OAI22_X1 U721 ( .A1(n2370), .A2(n1791), .B1(n2274), .B2(n1788), .ZN(n1547)
         );
  OAI22_X1 U722 ( .A1(n2306), .A2(n1779), .B1(n2402), .B2(n1776), .ZN(n1548)
         );
  OAI22_X1 U723 ( .A1(n2369), .A2(n1791), .B1(n2273), .B2(n1788), .ZN(n1564)
         );
  OAI22_X1 U724 ( .A1(n2305), .A2(n1779), .B1(n2401), .B2(n1776), .ZN(n1565)
         );
  OAI22_X1 U725 ( .A1(n2368), .A2(n1791), .B1(n2272), .B2(n1788), .ZN(n1581)
         );
  OAI22_X1 U726 ( .A1(n2304), .A2(n1779), .B1(n2400), .B2(n1776), .ZN(n1582)
         );
  OAI22_X1 U727 ( .A1(n2367), .A2(n1791), .B1(n2271), .B2(n1788), .ZN(n1598)
         );
  OAI22_X1 U728 ( .A1(n2303), .A2(n1779), .B1(n2399), .B2(n1776), .ZN(n1599)
         );
  OAI22_X1 U729 ( .A1(n2366), .A2(n1791), .B1(n2270), .B2(n1788), .ZN(n1615)
         );
  OAI22_X1 U730 ( .A1(n2302), .A2(n1779), .B1(n2398), .B2(n1776), .ZN(n1616)
         );
  OAI22_X1 U731 ( .A1(n2365), .A2(n1791), .B1(n2269), .B2(n1788), .ZN(n1632)
         );
  OAI22_X1 U732 ( .A1(n2301), .A2(n1779), .B1(n2397), .B2(n1776), .ZN(n1633)
         );
  OAI22_X1 U733 ( .A1(n2364), .A2(n1791), .B1(n2268), .B2(n1788), .ZN(n1649)
         );
  OAI22_X1 U734 ( .A1(n2300), .A2(n1779), .B1(n2396), .B2(n1776), .ZN(n1650)
         );
  OAI22_X1 U735 ( .A1(n2363), .A2(n1791), .B1(n2267), .B2(n1788), .ZN(n1666)
         );
  OAI22_X1 U736 ( .A1(n2299), .A2(n1779), .B1(n2395), .B2(n1776), .ZN(n1667)
         );
  OAI22_X1 U737 ( .A1(n2362), .A2(n1791), .B1(n2266), .B2(n1788), .ZN(n1683)
         );
  OAI22_X1 U738 ( .A1(n2298), .A2(n1779), .B1(n2394), .B2(n1776), .ZN(n1684)
         );
  OAI22_X1 U739 ( .A1(n2361), .A2(n1791), .B1(n2265), .B2(n1788), .ZN(n1711)
         );
  OAI22_X1 U740 ( .A1(n2297), .A2(n1779), .B1(n2393), .B2(n1776), .ZN(n1713)
         );
  OAI22_X1 U741 ( .A1(n1885), .A2(n2384), .B1(n1882), .B2(n2288), .ZN(n722) );
  OAI22_X1 U742 ( .A1(n1873), .A2(n2320), .B1(n1870), .B2(n2416), .ZN(n723) );
  OAI22_X1 U743 ( .A1(n1885), .A2(n2383), .B1(n1882), .B2(n2287), .ZN(n739) );
  OAI22_X1 U744 ( .A1(n1873), .A2(n2319), .B1(n1870), .B2(n2415), .ZN(n740) );
  OAI22_X1 U745 ( .A1(n1885), .A2(n2382), .B1(n1882), .B2(n2286), .ZN(n756) );
  OAI22_X1 U746 ( .A1(n1873), .A2(n2318), .B1(n1870), .B2(n2414), .ZN(n757) );
  OAI22_X1 U747 ( .A1(n1885), .A2(n2381), .B1(n1882), .B2(n2285), .ZN(n773) );
  OAI22_X1 U748 ( .A1(n1873), .A2(n2317), .B1(n1870), .B2(n2413), .ZN(n774) );
  OAI22_X1 U749 ( .A1(n1885), .A2(n2380), .B1(n1882), .B2(n2284), .ZN(n790) );
  OAI22_X1 U750 ( .A1(n1873), .A2(n2316), .B1(n1870), .B2(n2412), .ZN(n791) );
  OAI22_X1 U751 ( .A1(n1885), .A2(n2379), .B1(n1882), .B2(n2283), .ZN(n807) );
  OAI22_X1 U752 ( .A1(n1873), .A2(n2315), .B1(n1870), .B2(n2411), .ZN(n808) );
  OAI22_X1 U753 ( .A1(n1885), .A2(n2378), .B1(n1882), .B2(n2282), .ZN(n824) );
  OAI22_X1 U754 ( .A1(n1873), .A2(n2314), .B1(n1870), .B2(n2410), .ZN(n825) );
  OAI22_X1 U755 ( .A1(n1885), .A2(n2377), .B1(n1882), .B2(n2281), .ZN(n841) );
  OAI22_X1 U756 ( .A1(n1873), .A2(n2313), .B1(n1870), .B2(n2409), .ZN(n842) );
  OAI22_X1 U757 ( .A1(n1885), .A2(n2376), .B1(n1882), .B2(n2280), .ZN(n858) );
  OAI22_X1 U758 ( .A1(n1873), .A2(n2312), .B1(n1870), .B2(n2408), .ZN(n859) );
  OAI22_X1 U759 ( .A1(n1885), .A2(n2375), .B1(n1882), .B2(n2279), .ZN(n875) );
  OAI22_X1 U760 ( .A1(n1873), .A2(n2311), .B1(n1870), .B2(n2407), .ZN(n876) );
  OAI22_X1 U761 ( .A1(n1885), .A2(n2374), .B1(n1882), .B2(n2278), .ZN(n892) );
  OAI22_X1 U762 ( .A1(n1873), .A2(n2310), .B1(n1870), .B2(n2406), .ZN(n893) );
  OAI22_X1 U763 ( .A1(n1885), .A2(n2373), .B1(n1882), .B2(n2277), .ZN(n909) );
  OAI22_X1 U764 ( .A1(n1873), .A2(n2309), .B1(n1870), .B2(n2405), .ZN(n910) );
  OAI22_X1 U765 ( .A1(n1884), .A2(n2372), .B1(n1881), .B2(n2276), .ZN(n926) );
  OAI22_X1 U766 ( .A1(n1872), .A2(n2308), .B1(n1869), .B2(n2404), .ZN(n927) );
  OAI22_X1 U767 ( .A1(n1884), .A2(n2371), .B1(n1881), .B2(n2275), .ZN(n943) );
  OAI22_X1 U768 ( .A1(n1872), .A2(n2307), .B1(n1869), .B2(n2403), .ZN(n944) );
  OAI22_X1 U769 ( .A1(n1884), .A2(n2370), .B1(n1881), .B2(n2274), .ZN(n960) );
  OAI22_X1 U770 ( .A1(n1872), .A2(n2306), .B1(n1869), .B2(n2402), .ZN(n961) );
  OAI22_X1 U771 ( .A1(n1884), .A2(n2369), .B1(n1881), .B2(n2273), .ZN(n977) );
  OAI22_X1 U772 ( .A1(n1872), .A2(n2305), .B1(n1869), .B2(n2401), .ZN(n978) );
  OAI22_X1 U773 ( .A1(n1884), .A2(n2368), .B1(n1881), .B2(n2272), .ZN(n994) );
  OAI22_X1 U774 ( .A1(n1872), .A2(n2304), .B1(n1869), .B2(n2400), .ZN(n995) );
  OAI22_X1 U775 ( .A1(n1884), .A2(n2367), .B1(n1881), .B2(n2271), .ZN(n1011)
         );
  OAI22_X1 U776 ( .A1(n1872), .A2(n2303), .B1(n1869), .B2(n2399), .ZN(n1012)
         );
  OAI22_X1 U777 ( .A1(n1884), .A2(n2366), .B1(n1881), .B2(n2270), .ZN(n1028)
         );
  OAI22_X1 U778 ( .A1(n1872), .A2(n2302), .B1(n1869), .B2(n2398), .ZN(n1029)
         );
  OAI22_X1 U779 ( .A1(n1884), .A2(n2365), .B1(n1881), .B2(n2269), .ZN(n1045)
         );
  OAI22_X1 U780 ( .A1(n1872), .A2(n2301), .B1(n1869), .B2(n2397), .ZN(n1046)
         );
  OAI22_X1 U781 ( .A1(n1884), .A2(n2364), .B1(n1881), .B2(n2268), .ZN(n1062)
         );
  OAI22_X1 U782 ( .A1(n1872), .A2(n2300), .B1(n1869), .B2(n2396), .ZN(n1063)
         );
  OAI22_X1 U783 ( .A1(n1884), .A2(n2363), .B1(n1881), .B2(n2267), .ZN(n1079)
         );
  OAI22_X1 U784 ( .A1(n1872), .A2(n2299), .B1(n1869), .B2(n2395), .ZN(n1080)
         );
  OAI22_X1 U785 ( .A1(n1884), .A2(n2362), .B1(n1881), .B2(n2266), .ZN(n1096)
         );
  OAI22_X1 U786 ( .A1(n1872), .A2(n2298), .B1(n1869), .B2(n2394), .ZN(n1097)
         );
  OAI22_X1 U787 ( .A1(n1884), .A2(n2361), .B1(n1881), .B2(n2265), .ZN(n1124)
         );
  OAI22_X1 U788 ( .A1(n1872), .A2(n2297), .B1(n1869), .B2(n2393), .ZN(n1126)
         );
  OAI22_X1 U789 ( .A1(n2352), .A2(n1816), .B1(n2224), .B2(n1813), .ZN(n1307)
         );
  OAI22_X1 U790 ( .A1(n2351), .A2(n1816), .B1(n2223), .B2(n1813), .ZN(n1324)
         );
  OAI22_X1 U791 ( .A1(n2350), .A2(n1816), .B1(n2222), .B2(n1813), .ZN(n1341)
         );
  OAI22_X1 U792 ( .A1(n2349), .A2(n1816), .B1(n2221), .B2(n1813), .ZN(n1358)
         );
  OAI22_X1 U793 ( .A1(n2348), .A2(n1816), .B1(n2220), .B2(n1813), .ZN(n1375)
         );
  OAI22_X1 U794 ( .A1(n2347), .A2(n1816), .B1(n2219), .B2(n1813), .ZN(n1392)
         );
  OAI22_X1 U795 ( .A1(n2346), .A2(n1816), .B1(n2218), .B2(n1813), .ZN(n1409)
         );
  OAI22_X1 U796 ( .A1(n2345), .A2(n1816), .B1(n2217), .B2(n1813), .ZN(n1426)
         );
  OAI22_X1 U797 ( .A1(n2344), .A2(n1816), .B1(n2216), .B2(n1813), .ZN(n1443)
         );
  OAI22_X1 U798 ( .A1(n2343), .A2(n1816), .B1(n2215), .B2(n1813), .ZN(n1460)
         );
  OAI22_X1 U799 ( .A1(n2342), .A2(n1816), .B1(n2214), .B2(n1813), .ZN(n1477)
         );
  OAI22_X1 U800 ( .A1(n2341), .A2(n1816), .B1(n2213), .B2(n1813), .ZN(n1494)
         );
  OAI22_X1 U801 ( .A1(n2340), .A2(n1815), .B1(n2212), .B2(n1812), .ZN(n1511)
         );
  OAI22_X1 U802 ( .A1(n2339), .A2(n1815), .B1(n2211), .B2(n1812), .ZN(n1528)
         );
  OAI22_X1 U803 ( .A1(n2338), .A2(n1815), .B1(n2210), .B2(n1812), .ZN(n1545)
         );
  OAI22_X1 U804 ( .A1(n2337), .A2(n1815), .B1(n2209), .B2(n1812), .ZN(n1562)
         );
  OAI22_X1 U805 ( .A1(n2336), .A2(n1815), .B1(n2208), .B2(n1812), .ZN(n1579)
         );
  OAI22_X1 U806 ( .A1(n2335), .A2(n1815), .B1(n2207), .B2(n1812), .ZN(n1596)
         );
  OAI22_X1 U807 ( .A1(n2334), .A2(n1815), .B1(n2206), .B2(n1812), .ZN(n1613)
         );
  OAI22_X1 U808 ( .A1(n2333), .A2(n1815), .B1(n2205), .B2(n1812), .ZN(n1630)
         );
  OAI22_X1 U809 ( .A1(n2332), .A2(n1815), .B1(n2204), .B2(n1812), .ZN(n1647)
         );
  OAI22_X1 U810 ( .A1(n2331), .A2(n1815), .B1(n2203), .B2(n1812), .ZN(n1664)
         );
  OAI22_X1 U811 ( .A1(n2330), .A2(n1815), .B1(n2202), .B2(n1812), .ZN(n1681)
         );
  OAI22_X1 U812 ( .A1(n2329), .A2(n1815), .B1(n2201), .B2(n1812), .ZN(n1706)
         );
  OAI22_X1 U813 ( .A1(n1909), .A2(n2352), .B1(n1906), .B2(n2224), .ZN(n720) );
  OAI22_X1 U814 ( .A1(n1909), .A2(n2351), .B1(n1906), .B2(n2223), .ZN(n737) );
  OAI22_X1 U815 ( .A1(n1909), .A2(n2350), .B1(n1906), .B2(n2222), .ZN(n754) );
  OAI22_X1 U816 ( .A1(n1909), .A2(n2349), .B1(n1906), .B2(n2221), .ZN(n771) );
  OAI22_X1 U817 ( .A1(n1909), .A2(n2348), .B1(n1906), .B2(n2220), .ZN(n788) );
  OAI22_X1 U818 ( .A1(n1909), .A2(n2347), .B1(n1906), .B2(n2219), .ZN(n805) );
  OAI22_X1 U819 ( .A1(n1909), .A2(n2346), .B1(n1906), .B2(n2218), .ZN(n822) );
  OAI22_X1 U820 ( .A1(n1909), .A2(n2345), .B1(n1906), .B2(n2217), .ZN(n839) );
  OAI22_X1 U821 ( .A1(n1909), .A2(n2344), .B1(n1906), .B2(n2216), .ZN(n856) );
  OAI22_X1 U822 ( .A1(n1909), .A2(n2343), .B1(n1906), .B2(n2215), .ZN(n873) );
  OAI22_X1 U823 ( .A1(n1909), .A2(n2342), .B1(n1906), .B2(n2214), .ZN(n890) );
  OAI22_X1 U824 ( .A1(n1909), .A2(n2341), .B1(n1906), .B2(n2213), .ZN(n907) );
  OAI22_X1 U825 ( .A1(n1908), .A2(n2340), .B1(n1905), .B2(n2212), .ZN(n924) );
  OAI22_X1 U826 ( .A1(n1908), .A2(n2339), .B1(n1905), .B2(n2211), .ZN(n941) );
  OAI22_X1 U827 ( .A1(n1908), .A2(n2338), .B1(n1905), .B2(n2210), .ZN(n958) );
  OAI22_X1 U828 ( .A1(n1908), .A2(n2337), .B1(n1905), .B2(n2209), .ZN(n975) );
  OAI22_X1 U829 ( .A1(n1908), .A2(n2336), .B1(n1905), .B2(n2208), .ZN(n992) );
  OAI22_X1 U830 ( .A1(n1908), .A2(n2335), .B1(n1905), .B2(n2207), .ZN(n1009)
         );
  OAI22_X1 U831 ( .A1(n1908), .A2(n2334), .B1(n1905), .B2(n2206), .ZN(n1026)
         );
  OAI22_X1 U832 ( .A1(n1908), .A2(n2333), .B1(n1905), .B2(n2205), .ZN(n1043)
         );
  OAI22_X1 U833 ( .A1(n1908), .A2(n2332), .B1(n1905), .B2(n2204), .ZN(n1060)
         );
  OAI22_X1 U834 ( .A1(n1908), .A2(n2331), .B1(n1905), .B2(n2203), .ZN(n1077)
         );
  OAI22_X1 U835 ( .A1(n1908), .A2(n2330), .B1(n1905), .B2(n2202), .ZN(n1094)
         );
  OAI22_X1 U836 ( .A1(n1908), .A2(n2329), .B1(n1905), .B2(n2201), .ZN(n1119)
         );
  NAND2_X1 U837 ( .A1(n1697), .A2(n1702), .ZN(n1146) );
  NAND2_X1 U838 ( .A1(n1697), .A2(n1703), .ZN(n1145) );
  NAND2_X1 U839 ( .A1(n1110), .A2(n1116), .ZN(n558) );
  NAND2_X1 U840 ( .A1(n1110), .A2(n1115), .ZN(n559) );
  NAND2_X1 U841 ( .A1(n1700), .A2(n1703), .ZN(n1150) );
  NAND2_X1 U842 ( .A1(n1113), .A2(n1116), .ZN(n563) );
  NAND2_X1 U843 ( .A1(n1708), .A2(n1695), .ZN(n1169) );
  NAND2_X1 U844 ( .A1(n1708), .A2(n1699), .ZN(n1174) );
  NAND2_X1 U845 ( .A1(n1708), .A2(n1697), .ZN(n1158) );
  NAND2_X1 U846 ( .A1(n1121), .A2(n1108), .ZN(n582) );
  NAND2_X1 U847 ( .A1(n1121), .A2(n1112), .ZN(n587) );
  NAND2_X1 U848 ( .A1(n1121), .A2(n1110), .ZN(n571) );
  NAND2_X1 U849 ( .A1(n1712), .A2(n1697), .ZN(n1168) );
  NAND2_X1 U850 ( .A1(n1712), .A2(n1695), .ZN(n1173) );
  NAND2_X1 U851 ( .A1(n1710), .A2(n1699), .ZN(n1161) );
  NAND2_X1 U852 ( .A1(n1710), .A2(n1695), .ZN(n1160) );
  NAND2_X1 U853 ( .A1(n1125), .A2(n1110), .ZN(n581) );
  NAND2_X1 U854 ( .A1(n1125), .A2(n1108), .ZN(n586) );
  NAND2_X1 U855 ( .A1(n1123), .A2(n1108), .ZN(n573) );
  NAND2_X1 U856 ( .A1(n1123), .A2(n1112), .ZN(n574) );
  NAND2_X1 U857 ( .A1(n1694), .A2(n1697), .ZN(n1136) );
  NAND2_X1 U858 ( .A1(n1696), .A2(n1697), .ZN(n1135) );
  NAND2_X1 U859 ( .A1(n1109), .A2(n1110), .ZN(n548) );
  NAND2_X1 U860 ( .A1(n1107), .A2(n1110), .ZN(n549) );
  NAND2_X1 U861 ( .A1(n1707), .A2(n1700), .ZN(n1159) );
  NAND2_X1 U862 ( .A1(n1694), .A2(n1700), .ZN(n1141) );
  NAND2_X1 U863 ( .A1(n1696), .A2(n1700), .ZN(n1140) );
  NAND2_X1 U864 ( .A1(n1702), .A2(n1700), .ZN(n1151) );
  NAND2_X1 U865 ( .A1(n1109), .A2(n1113), .ZN(n553) );
  NAND2_X1 U866 ( .A1(n1107), .A2(n1113), .ZN(n554) );
  NAND2_X1 U867 ( .A1(n1115), .A2(n1113), .ZN(n564) );
  NAND2_X1 U868 ( .A1(n1120), .A2(n1113), .ZN(n572) );
  AND2_X1 U869 ( .A1(n1708), .A2(n1700), .ZN(n1166) );
  AND2_X1 U870 ( .A1(n1121), .A2(n1113), .ZN(n579) );
  AND2_X1 U871 ( .A1(n1699), .A2(n1703), .ZN(n1153) );
  AND2_X1 U872 ( .A1(n1699), .A2(n1702), .ZN(n1154) );
  AND2_X1 U873 ( .A1(n1112), .A2(n1116), .ZN(n566) );
  AND2_X1 U874 ( .A1(n1112), .A2(n1115), .ZN(n567) );
  AND2_X1 U875 ( .A1(n1710), .A2(n1697), .ZN(n1163) );
  AND2_X1 U876 ( .A1(n1712), .A2(n1699), .ZN(n1165) );
  AND2_X1 U877 ( .A1(n1712), .A2(n1700), .ZN(n1170) );
  AND2_X1 U878 ( .A1(n1710), .A2(n1700), .ZN(n1155) );
  AND2_X1 U879 ( .A1(n1108), .A2(n1116), .ZN(n561) );
  AND2_X1 U880 ( .A1(n1108), .A2(n1115), .ZN(n562) );
  AND2_X1 U881 ( .A1(n1695), .A2(n1703), .ZN(n1148) );
  AND2_X1 U882 ( .A1(n1695), .A2(n1702), .ZN(n1149) );
  AND2_X1 U883 ( .A1(n1123), .A2(n1110), .ZN(n576) );
  AND2_X1 U884 ( .A1(n1707), .A2(n1697), .ZN(n1171) );
  AND2_X1 U885 ( .A1(n1120), .A2(n1110), .ZN(n584) );
  AND2_X1 U886 ( .A1(n1125), .A2(n1112), .ZN(n578) );
  AND2_X1 U887 ( .A1(n1125), .A2(n1113), .ZN(n583) );
  AND2_X1 U888 ( .A1(n1123), .A2(n1113), .ZN(n568) );
  AND2_X1 U889 ( .A1(n1696), .A2(n1699), .ZN(n1143) );
  AND2_X1 U890 ( .A1(n1694), .A2(n1699), .ZN(n1144) );
  AND2_X1 U891 ( .A1(n1707), .A2(n1699), .ZN(n1164) );
  AND2_X1 U892 ( .A1(n1109), .A2(n1112), .ZN(n556) );
  AND2_X1 U893 ( .A1(n1107), .A2(n1112), .ZN(n557) );
  AND2_X1 U894 ( .A1(n1120), .A2(n1112), .ZN(n577) );
  AND2_X1 U895 ( .A1(n1109), .A2(n1108), .ZN(n551) );
  AND2_X1 U896 ( .A1(n1107), .A2(n1108), .ZN(n552) );
  AND2_X1 U897 ( .A1(n1696), .A2(n1695), .ZN(n1138) );
  AND2_X1 U898 ( .A1(n1694), .A2(n1695), .ZN(n1139) );
  OAI21_X1 U899 ( .B1(n533), .B2(n539), .A(n2161), .ZN(N340) );
  OAI21_X1 U900 ( .B1(n532), .B2(n539), .A(n2161), .ZN(N341) );
  OAI21_X1 U901 ( .B1(n531), .B2(n539), .A(n2161), .ZN(N342) );
  OAI21_X1 U902 ( .B1(n530), .B2(n539), .A(n2161), .ZN(N343) );
  OAI21_X1 U903 ( .B1(n529), .B2(n539), .A(n2161), .ZN(N344) );
  OAI21_X1 U904 ( .B1(n528), .B2(n539), .A(n2161), .ZN(N345) );
  OAI21_X1 U905 ( .B1(n534), .B2(n538), .A(n2161), .ZN(N347) );
  OAI21_X1 U906 ( .B1(n534), .B2(n539), .A(n2159), .ZN(N307) );
  OAI21_X1 U907 ( .B1(n537), .B2(n539), .A(n2160), .ZN(N346) );
  OAI21_X1 U908 ( .B1(n533), .B2(n538), .A(n2160), .ZN(N348) );
  OAI21_X1 U909 ( .B1(n532), .B2(n538), .A(n2160), .ZN(N349) );
  OAI21_X1 U910 ( .B1(n531), .B2(n538), .A(n2160), .ZN(N350) );
  OAI21_X1 U911 ( .B1(n530), .B2(n538), .A(n2160), .ZN(N351) );
  OAI21_X1 U912 ( .B1(n529), .B2(n538), .A(n2160), .ZN(N352) );
  OAI21_X1 U913 ( .B1(n528), .B2(n538), .A(n2160), .ZN(N353) );
  OAI21_X1 U914 ( .B1(n537), .B2(n538), .A(n2160), .ZN(N354) );
  OAI21_X1 U915 ( .B1(n534), .B2(n536), .A(n2160), .ZN(N355) );
  OAI21_X1 U916 ( .B1(n533), .B2(n536), .A(n2160), .ZN(N356) );
  OAI21_X1 U917 ( .B1(n532), .B2(n536), .A(n2160), .ZN(N357) );
  OAI21_X1 U918 ( .B1(n531), .B2(n536), .A(n2159), .ZN(N358) );
  OAI21_X1 U919 ( .B1(n530), .B2(n536), .A(n2160), .ZN(N359) );
  OAI21_X1 U920 ( .B1(n529), .B2(n536), .A(n2159), .ZN(N360) );
  OAI21_X1 U921 ( .B1(n528), .B2(n536), .A(n2159), .ZN(N361) );
  OAI21_X1 U922 ( .B1(n536), .B2(n537), .A(n2159), .ZN(N362) );
  OAI21_X1 U923 ( .B1(n527), .B2(n534), .A(n2159), .ZN(N363) );
  OAI21_X1 U924 ( .B1(n527), .B2(n533), .A(n2159), .ZN(N364) );
  OAI21_X1 U925 ( .B1(n527), .B2(n532), .A(n2159), .ZN(N365) );
  OAI21_X1 U926 ( .B1(n527), .B2(n531), .A(n2159), .ZN(N366) );
  OAI21_X1 U927 ( .B1(n527), .B2(n530), .A(n2159), .ZN(N367) );
  OAI21_X1 U928 ( .B1(n527), .B2(n529), .A(n2159), .ZN(N368) );
  OAI21_X1 U929 ( .B1(n527), .B2(n528), .A(n2159), .ZN(N369) );
  AND2_X1 U930 ( .A1(n2689), .A2(n2162), .ZN(N371) );
  AND2_X1 U931 ( .A1(datain[0]), .A2(n2161), .ZN(N308) );
  AND2_X1 U932 ( .A1(datain[15]), .A2(n2161), .ZN(N323) );
  AND2_X1 U933 ( .A1(datain[26]), .A2(n2161), .ZN(N334) );
  AND2_X1 U934 ( .A1(datain[27]), .A2(n2161), .ZN(N335) );
  AND2_X1 U935 ( .A1(datain[28]), .A2(n2161), .ZN(N336) );
  AND2_X1 U936 ( .A1(datain[29]), .A2(n2161), .ZN(N337) );
  AND2_X1 U937 ( .A1(datain[30]), .A2(n2161), .ZN(N338) );
  AND2_X1 U938 ( .A1(datain[31]), .A2(n2161), .ZN(N339) );
  AND2_X1 U939 ( .A1(datain[8]), .A2(n2162), .ZN(N316) );
  AND2_X1 U940 ( .A1(datain[9]), .A2(n2162), .ZN(N317) );
  AND2_X1 U941 ( .A1(datain[10]), .A2(n2162), .ZN(N318) );
  AND2_X1 U942 ( .A1(datain[11]), .A2(n2162), .ZN(N319) );
  AND2_X1 U943 ( .A1(datain[12]), .A2(n2162), .ZN(N320) );
  AND2_X1 U944 ( .A1(datain[13]), .A2(n2162), .ZN(N321) );
  AND2_X1 U945 ( .A1(datain[14]), .A2(n2162), .ZN(N322) );
  AND2_X1 U946 ( .A1(datain[16]), .A2(n2162), .ZN(N324) );
  AND2_X1 U947 ( .A1(datain[17]), .A2(n2162), .ZN(N325) );
  AND2_X1 U948 ( .A1(datain[18]), .A2(n2162), .ZN(N326) );
  AND2_X1 U949 ( .A1(datain[19]), .A2(n2162), .ZN(N327) );
  AND2_X1 U950 ( .A1(datain[20]), .A2(n2162), .ZN(N328) );
  AND2_X1 U951 ( .A1(datain[21]), .A2(n2162), .ZN(N329) );
  AND2_X1 U952 ( .A1(datain[22]), .A2(n2162), .ZN(N330) );
  AND2_X1 U953 ( .A1(datain[23]), .A2(n2162), .ZN(N331) );
  AND2_X1 U954 ( .A1(datain[24]), .A2(n2162), .ZN(N332) );
  AND2_X1 U955 ( .A1(datain[25]), .A2(n2162), .ZN(N333) );
  AND2_X1 U956 ( .A1(datain[1]), .A2(n2163), .ZN(N309) );
  AND2_X1 U957 ( .A1(datain[2]), .A2(n2163), .ZN(N310) );
  AND2_X1 U958 ( .A1(datain[3]), .A2(n2163), .ZN(N311) );
  AND2_X1 U959 ( .A1(datain[4]), .A2(n2163), .ZN(N312) );
  AND2_X1 U960 ( .A1(datain[5]), .A2(n2163), .ZN(N313) );
  AND2_X1 U961 ( .A1(datain[6]), .A2(n2163), .ZN(N314) );
  AND2_X1 U962 ( .A1(datain[7]), .A2(n2163), .ZN(N315) );
  NOR2_X1 U963 ( .A1(n2682), .A2(add_rd1[1]), .ZN(n1700) );
  NOR2_X1 U964 ( .A1(n2686), .A2(add_rd2[1]), .ZN(n1113) );
  NOR3_X1 U965 ( .A1(add_rd1[0]), .A2(add_rd1[4]), .A3(n2681), .ZN(n1708) );
  NOR3_X1 U966 ( .A1(add_rd2[0]), .A2(add_rd2[4]), .A3(n2685), .ZN(n1121) );
  NOR3_X1 U967 ( .A1(add_rd1[3]), .A2(add_rd1[4]), .A3(n2684), .ZN(n1710) );
  NOR3_X1 U968 ( .A1(n2684), .A2(add_rd1[4]), .A3(n2681), .ZN(n1712) );
  NOR2_X1 U969 ( .A1(add_rd2[1]), .A2(add_rd2[2]), .ZN(n1108) );
  NOR2_X1 U970 ( .A1(add_rd1[1]), .A2(add_rd1[2]), .ZN(n1695) );
  NOR3_X1 U971 ( .A1(add_rd2[3]), .A2(add_rd2[4]), .A3(n2688), .ZN(n1123) );
  NOR3_X1 U972 ( .A1(n2688), .A2(add_rd2[4]), .A3(n2685), .ZN(n1125) );
  NOR3_X1 U973 ( .A1(add_rd1[3]), .A2(add_rd1[4]), .A3(add_rd1[0]), .ZN(n1707)
         );
  NOR3_X1 U974 ( .A1(add_rd2[3]), .A2(add_rd2[4]), .A3(add_rd2[0]), .ZN(n1120)
         );
  OAI221_X1 U975 ( .B1(n1961), .B2(n2488), .C1(n1958), .C2(n2456), .A(n550), 
        .ZN(n547) );
  AOI22_X1 U976 ( .A1(\registers[17][0] ), .A2(n1955), .B1(\registers[16][0] ), 
        .B2(n1952), .ZN(n550) );
  OAI221_X1 U977 ( .B1(n1961), .B2(n2487), .C1(n1958), .C2(n2455), .A(n596), 
        .ZN(n595) );
  AOI22_X1 U978 ( .A1(\registers[17][1] ), .A2(n1955), .B1(\registers[16][1] ), 
        .B2(n1952), .ZN(n596) );
  OAI221_X1 U979 ( .B1(n1961), .B2(n2486), .C1(n1958), .C2(n2454), .A(n613), 
        .ZN(n612) );
  AOI22_X1 U980 ( .A1(\registers[17][2] ), .A2(n1955), .B1(\registers[16][2] ), 
        .B2(n1952), .ZN(n613) );
  OAI221_X1 U981 ( .B1(n1961), .B2(n2485), .C1(n1958), .C2(n2453), .A(n630), 
        .ZN(n629) );
  AOI22_X1 U982 ( .A1(\registers[17][3] ), .A2(n1955), .B1(\registers[16][3] ), 
        .B2(n1952), .ZN(n630) );
  OAI221_X1 U983 ( .B1(n1961), .B2(n2484), .C1(n1958), .C2(n2452), .A(n647), 
        .ZN(n646) );
  AOI22_X1 U984 ( .A1(\registers[17][4] ), .A2(n1955), .B1(\registers[16][4] ), 
        .B2(n1952), .ZN(n647) );
  OAI221_X1 U985 ( .B1(n1961), .B2(n2483), .C1(n1958), .C2(n2451), .A(n664), 
        .ZN(n663) );
  AOI22_X1 U986 ( .A1(\registers[17][5] ), .A2(n1955), .B1(\registers[16][5] ), 
        .B2(n1952), .ZN(n664) );
  OAI221_X1 U987 ( .B1(n1961), .B2(n2482), .C1(n1958), .C2(n2450), .A(n681), 
        .ZN(n680) );
  AOI22_X1 U988 ( .A1(\registers[17][6] ), .A2(n1955), .B1(\registers[16][6] ), 
        .B2(n1952), .ZN(n681) );
  OAI221_X1 U989 ( .B1(n1961), .B2(n2481), .C1(n1958), .C2(n2449), .A(n698), 
        .ZN(n697) );
  AOI22_X1 U990 ( .A1(\registers[17][7] ), .A2(n1955), .B1(\registers[16][7] ), 
        .B2(n1952), .ZN(n698) );
  OAI221_X1 U991 ( .B1(n2488), .B2(n1868), .C1(n2456), .C2(n1865), .A(n1137), 
        .ZN(n1134) );
  AOI22_X1 U992 ( .A1(n1862), .A2(\registers[17][0] ), .B1(n1857), .B2(
        \registers[16][0] ), .ZN(n1137) );
  OAI221_X1 U993 ( .B1(n2487), .B2(n1868), .C1(n2455), .C2(n1865), .A(n1183), 
        .ZN(n1182) );
  AOI22_X1 U994 ( .A1(n1862), .A2(\registers[17][1] ), .B1(n1857), .B2(
        \registers[16][1] ), .ZN(n1183) );
  OAI221_X1 U995 ( .B1(n2486), .B2(n1868), .C1(n2454), .C2(n1865), .A(n1200), 
        .ZN(n1199) );
  AOI22_X1 U996 ( .A1(n1862), .A2(\registers[17][2] ), .B1(n1857), .B2(
        \registers[16][2] ), .ZN(n1200) );
  OAI221_X1 U997 ( .B1(n2485), .B2(n1868), .C1(n2453), .C2(n1865), .A(n1217), 
        .ZN(n1216) );
  AOI22_X1 U998 ( .A1(n1862), .A2(\registers[17][3] ), .B1(n1857), .B2(
        \registers[16][3] ), .ZN(n1217) );
  OAI221_X1 U999 ( .B1(n2484), .B2(n1868), .C1(n2452), .C2(n1865), .A(n1234), 
        .ZN(n1233) );
  AOI22_X1 U1000 ( .A1(n1862), .A2(\registers[17][4] ), .B1(n1857), .B2(
        \registers[16][4] ), .ZN(n1234) );
  OAI221_X1 U1001 ( .B1(n2483), .B2(n1868), .C1(n2451), .C2(n1865), .A(n1251), 
        .ZN(n1250) );
  AOI22_X1 U1002 ( .A1(n1862), .A2(\registers[17][5] ), .B1(n1857), .B2(
        \registers[16][5] ), .ZN(n1251) );
  OAI221_X1 U1003 ( .B1(n2482), .B2(n1868), .C1(n2450), .C2(n1865), .A(n1268), 
        .ZN(n1267) );
  AOI22_X1 U1004 ( .A1(n1862), .A2(\registers[17][6] ), .B1(n1857), .B2(
        \registers[16][6] ), .ZN(n1268) );
  OAI221_X1 U1005 ( .B1(n2481), .B2(n1868), .C1(n2449), .C2(n1865), .A(n1285), 
        .ZN(n1284) );
  AOI22_X1 U1006 ( .A1(n1862), .A2(\registers[17][7] ), .B1(n1857), .B2(
        \registers[16][7] ), .ZN(n1285) );
  OAI221_X1 U1007 ( .B1(n2480), .B2(n1867), .C1(n2448), .C2(n1864), .A(n1302), 
        .ZN(n1301) );
  AOI22_X1 U1008 ( .A1(n1861), .A2(\registers[17][8] ), .B1(n1857), .B2(
        \registers[16][8] ), .ZN(n1302) );
  OAI221_X1 U1009 ( .B1(n2479), .B2(n1867), .C1(n2447), .C2(n1864), .A(n1319), 
        .ZN(n1318) );
  AOI22_X1 U1010 ( .A1(n1861), .A2(\registers[17][9] ), .B1(n1857), .B2(
        \registers[16][9] ), .ZN(n1319) );
  OAI221_X1 U1011 ( .B1(n2478), .B2(n1867), .C1(n2446), .C2(n1864), .A(n1336), 
        .ZN(n1335) );
  AOI22_X1 U1012 ( .A1(n1861), .A2(\registers[17][10] ), .B1(n1857), .B2(
        \registers[16][10] ), .ZN(n1336) );
  OAI221_X1 U1013 ( .B1(n2477), .B2(n1867), .C1(n2445), .C2(n1864), .A(n1353), 
        .ZN(n1352) );
  AOI22_X1 U1014 ( .A1(n1861), .A2(\registers[17][11] ), .B1(n1857), .B2(
        \registers[16][11] ), .ZN(n1353) );
  OAI221_X1 U1015 ( .B1(n2476), .B2(n1867), .C1(n2444), .C2(n1864), .A(n1370), 
        .ZN(n1369) );
  AOI22_X1 U1016 ( .A1(n1861), .A2(\registers[17][12] ), .B1(n1858), .B2(
        \registers[16][12] ), .ZN(n1370) );
  OAI221_X1 U1017 ( .B1(n2475), .B2(n1867), .C1(n2443), .C2(n1864), .A(n1387), 
        .ZN(n1386) );
  AOI22_X1 U1018 ( .A1(n1861), .A2(\registers[17][13] ), .B1(n1858), .B2(
        \registers[16][13] ), .ZN(n1387) );
  OAI221_X1 U1019 ( .B1(n2474), .B2(n1867), .C1(n2442), .C2(n1864), .A(n1404), 
        .ZN(n1403) );
  AOI22_X1 U1020 ( .A1(n1861), .A2(\registers[17][14] ), .B1(n1858), .B2(
        \registers[16][14] ), .ZN(n1404) );
  OAI221_X1 U1021 ( .B1(n2473), .B2(n1867), .C1(n2441), .C2(n1864), .A(n1421), 
        .ZN(n1420) );
  AOI22_X1 U1022 ( .A1(n1861), .A2(\registers[17][15] ), .B1(n1858), .B2(
        \registers[16][15] ), .ZN(n1421) );
  OAI221_X1 U1023 ( .B1(n2472), .B2(n1867), .C1(n2440), .C2(n1864), .A(n1438), 
        .ZN(n1437) );
  AOI22_X1 U1024 ( .A1(n1861), .A2(\registers[17][16] ), .B1(n1858), .B2(
        \registers[16][16] ), .ZN(n1438) );
  OAI221_X1 U1025 ( .B1(n2471), .B2(n1867), .C1(n2439), .C2(n1864), .A(n1455), 
        .ZN(n1454) );
  AOI22_X1 U1026 ( .A1(n1861), .A2(\registers[17][17] ), .B1(n1858), .B2(
        \registers[16][17] ), .ZN(n1455) );
  OAI221_X1 U1027 ( .B1(n2470), .B2(n1867), .C1(n2438), .C2(n1864), .A(n1472), 
        .ZN(n1471) );
  AOI22_X1 U1028 ( .A1(n1861), .A2(\registers[17][18] ), .B1(n1858), .B2(
        \registers[16][18] ), .ZN(n1472) );
  OAI221_X1 U1029 ( .B1(n2469), .B2(n1867), .C1(n2437), .C2(n1864), .A(n1489), 
        .ZN(n1488) );
  AOI22_X1 U1030 ( .A1(n1861), .A2(\registers[17][19] ), .B1(n1858), .B2(
        \registers[16][19] ), .ZN(n1489) );
  OAI221_X1 U1031 ( .B1(n2468), .B2(n1866), .C1(n2436), .C2(n1863), .A(n1506), 
        .ZN(n1505) );
  AOI22_X1 U1032 ( .A1(n1860), .A2(\registers[17][20] ), .B1(n1858), .B2(
        \registers[16][20] ), .ZN(n1506) );
  OAI221_X1 U1033 ( .B1(n2467), .B2(n1866), .C1(n2435), .C2(n1863), .A(n1523), 
        .ZN(n1522) );
  AOI22_X1 U1034 ( .A1(n1860), .A2(\registers[17][21] ), .B1(n1858), .B2(
        \registers[16][21] ), .ZN(n1523) );
  OAI221_X1 U1035 ( .B1(n2466), .B2(n1866), .C1(n2434), .C2(n1863), .A(n1540), 
        .ZN(n1539) );
  AOI22_X1 U1036 ( .A1(n1860), .A2(\registers[17][22] ), .B1(n1858), .B2(
        \registers[16][22] ), .ZN(n1540) );
  OAI221_X1 U1037 ( .B1(n2465), .B2(n1866), .C1(n2433), .C2(n1863), .A(n1557), 
        .ZN(n1556) );
  AOI22_X1 U1038 ( .A1(n1860), .A2(\registers[17][23] ), .B1(n1858), .B2(
        \registers[16][23] ), .ZN(n1557) );
  OAI221_X1 U1039 ( .B1(n2464), .B2(n1866), .C1(n2432), .C2(n1863), .A(n1574), 
        .ZN(n1573) );
  AOI22_X1 U1040 ( .A1(n1860), .A2(\registers[17][24] ), .B1(n1859), .B2(
        \registers[16][24] ), .ZN(n1574) );
  OAI221_X1 U1041 ( .B1(n2463), .B2(n1866), .C1(n2431), .C2(n1863), .A(n1591), 
        .ZN(n1590) );
  AOI22_X1 U1042 ( .A1(n1860), .A2(\registers[17][25] ), .B1(n1859), .B2(
        \registers[16][25] ), .ZN(n1591) );
  OAI221_X1 U1043 ( .B1(n2462), .B2(n1866), .C1(n2430), .C2(n1863), .A(n1608), 
        .ZN(n1607) );
  AOI22_X1 U1044 ( .A1(n1860), .A2(\registers[17][26] ), .B1(n1859), .B2(
        \registers[16][26] ), .ZN(n1608) );
  OAI221_X1 U1045 ( .B1(n2461), .B2(n1866), .C1(n2429), .C2(n1863), .A(n1625), 
        .ZN(n1624) );
  AOI22_X1 U1046 ( .A1(n1860), .A2(\registers[17][27] ), .B1(n1859), .B2(
        \registers[16][27] ), .ZN(n1625) );
  OAI221_X1 U1047 ( .B1(n2460), .B2(n1866), .C1(n2428), .C2(n1863), .A(n1642), 
        .ZN(n1641) );
  AOI22_X1 U1048 ( .A1(n1860), .A2(\registers[17][28] ), .B1(n1859), .B2(
        \registers[16][28] ), .ZN(n1642) );
  OAI221_X1 U1049 ( .B1(n2459), .B2(n1866), .C1(n2427), .C2(n1863), .A(n1659), 
        .ZN(n1658) );
  AOI22_X1 U1050 ( .A1(n1860), .A2(\registers[17][29] ), .B1(n1859), .B2(
        \registers[16][29] ), .ZN(n1659) );
  OAI221_X1 U1051 ( .B1(n2458), .B2(n1866), .C1(n2426), .C2(n1863), .A(n1676), 
        .ZN(n1675) );
  AOI22_X1 U1052 ( .A1(n1860), .A2(\registers[17][30] ), .B1(n1859), .B2(
        \registers[16][30] ), .ZN(n1676) );
  OAI221_X1 U1053 ( .B1(n2457), .B2(n1866), .C1(n2425), .C2(n1863), .A(n1693), 
        .ZN(n1692) );
  AOI22_X1 U1054 ( .A1(n1860), .A2(\registers[17][31] ), .B1(n1859), .B2(
        \registers[16][31] ), .ZN(n1693) );
  OAI221_X1 U1055 ( .B1(n1960), .B2(n2480), .C1(n1957), .C2(n2448), .A(n715), 
        .ZN(n714) );
  AOI22_X1 U1056 ( .A1(\registers[17][8] ), .A2(n1954), .B1(\registers[16][8] ), .B2(n1951), .ZN(n715) );
  OAI221_X1 U1057 ( .B1(n1960), .B2(n2479), .C1(n1957), .C2(n2447), .A(n732), 
        .ZN(n731) );
  AOI22_X1 U1058 ( .A1(\registers[17][9] ), .A2(n1954), .B1(\registers[16][9] ), .B2(n1951), .ZN(n732) );
  OAI221_X1 U1059 ( .B1(n1960), .B2(n2478), .C1(n1957), .C2(n2446), .A(n749), 
        .ZN(n748) );
  AOI22_X1 U1060 ( .A1(\registers[17][10] ), .A2(n1954), .B1(
        \registers[16][10] ), .B2(n1951), .ZN(n749) );
  OAI221_X1 U1061 ( .B1(n1960), .B2(n2477), .C1(n1957), .C2(n2445), .A(n766), 
        .ZN(n765) );
  AOI22_X1 U1062 ( .A1(\registers[17][11] ), .A2(n1954), .B1(
        \registers[16][11] ), .B2(n1951), .ZN(n766) );
  OAI221_X1 U1063 ( .B1(n1960), .B2(n2476), .C1(n1957), .C2(n2444), .A(n783), 
        .ZN(n782) );
  AOI22_X1 U1064 ( .A1(\registers[17][12] ), .A2(n1954), .B1(
        \registers[16][12] ), .B2(n1951), .ZN(n783) );
  OAI221_X1 U1065 ( .B1(n1960), .B2(n2475), .C1(n1957), .C2(n2443), .A(n800), 
        .ZN(n799) );
  AOI22_X1 U1066 ( .A1(\registers[17][13] ), .A2(n1954), .B1(
        \registers[16][13] ), .B2(n1951), .ZN(n800) );
  OAI221_X1 U1067 ( .B1(n1960), .B2(n2474), .C1(n1957), .C2(n2442), .A(n817), 
        .ZN(n816) );
  AOI22_X1 U1068 ( .A1(\registers[17][14] ), .A2(n1954), .B1(
        \registers[16][14] ), .B2(n1951), .ZN(n817) );
  OAI221_X1 U1069 ( .B1(n1960), .B2(n2473), .C1(n1957), .C2(n2441), .A(n834), 
        .ZN(n833) );
  AOI22_X1 U1070 ( .A1(\registers[17][15] ), .A2(n1954), .B1(
        \registers[16][15] ), .B2(n1951), .ZN(n834) );
  OAI221_X1 U1071 ( .B1(n1960), .B2(n2472), .C1(n1957), .C2(n2440), .A(n851), 
        .ZN(n850) );
  AOI22_X1 U1072 ( .A1(\registers[17][16] ), .A2(n1954), .B1(
        \registers[16][16] ), .B2(n1951), .ZN(n851) );
  OAI221_X1 U1073 ( .B1(n1960), .B2(n2471), .C1(n1957), .C2(n2439), .A(n868), 
        .ZN(n867) );
  AOI22_X1 U1074 ( .A1(\registers[17][17] ), .A2(n1954), .B1(
        \registers[16][17] ), .B2(n1951), .ZN(n868) );
  OAI221_X1 U1075 ( .B1(n1960), .B2(n2470), .C1(n1957), .C2(n2438), .A(n885), 
        .ZN(n884) );
  AOI22_X1 U1076 ( .A1(\registers[17][18] ), .A2(n1954), .B1(
        \registers[16][18] ), .B2(n1951), .ZN(n885) );
  OAI221_X1 U1077 ( .B1(n1960), .B2(n2469), .C1(n1957), .C2(n2437), .A(n902), 
        .ZN(n901) );
  AOI22_X1 U1078 ( .A1(\registers[17][19] ), .A2(n1954), .B1(
        \registers[16][19] ), .B2(n1951), .ZN(n902) );
  OAI221_X1 U1079 ( .B1(n1959), .B2(n2468), .C1(n1956), .C2(n2436), .A(n919), 
        .ZN(n918) );
  AOI22_X1 U1080 ( .A1(\registers[17][20] ), .A2(n1953), .B1(
        \registers[16][20] ), .B2(n1950), .ZN(n919) );
  OAI221_X1 U1081 ( .B1(n1959), .B2(n2467), .C1(n1956), .C2(n2435), .A(n936), 
        .ZN(n935) );
  AOI22_X1 U1082 ( .A1(\registers[17][21] ), .A2(n1953), .B1(
        \registers[16][21] ), .B2(n1950), .ZN(n936) );
  OAI221_X1 U1083 ( .B1(n1959), .B2(n2466), .C1(n1956), .C2(n2434), .A(n953), 
        .ZN(n952) );
  AOI22_X1 U1084 ( .A1(\registers[17][22] ), .A2(n1953), .B1(
        \registers[16][22] ), .B2(n1950), .ZN(n953) );
  OAI221_X1 U1085 ( .B1(n1959), .B2(n2465), .C1(n1956), .C2(n2433), .A(n970), 
        .ZN(n969) );
  AOI22_X1 U1086 ( .A1(\registers[17][23] ), .A2(n1953), .B1(
        \registers[16][23] ), .B2(n1950), .ZN(n970) );
  OAI221_X1 U1087 ( .B1(n1959), .B2(n2464), .C1(n1956), .C2(n2432), .A(n987), 
        .ZN(n986) );
  AOI22_X1 U1088 ( .A1(\registers[17][24] ), .A2(n1953), .B1(
        \registers[16][24] ), .B2(n1950), .ZN(n987) );
  OAI221_X1 U1089 ( .B1(n1959), .B2(n2463), .C1(n1956), .C2(n2431), .A(n1004), 
        .ZN(n1003) );
  AOI22_X1 U1090 ( .A1(\registers[17][25] ), .A2(n1953), .B1(
        \registers[16][25] ), .B2(n1950), .ZN(n1004) );
  OAI221_X1 U1091 ( .B1(n1959), .B2(n2462), .C1(n1956), .C2(n2430), .A(n1021), 
        .ZN(n1020) );
  AOI22_X1 U1092 ( .A1(\registers[17][26] ), .A2(n1953), .B1(
        \registers[16][26] ), .B2(n1950), .ZN(n1021) );
  OAI221_X1 U1093 ( .B1(n1959), .B2(n2461), .C1(n1956), .C2(n2429), .A(n1038), 
        .ZN(n1037) );
  AOI22_X1 U1094 ( .A1(\registers[17][27] ), .A2(n1953), .B1(
        \registers[16][27] ), .B2(n1950), .ZN(n1038) );
  OAI221_X1 U1095 ( .B1(n1959), .B2(n2460), .C1(n1956), .C2(n2428), .A(n1055), 
        .ZN(n1054) );
  AOI22_X1 U1096 ( .A1(\registers[17][28] ), .A2(n1953), .B1(
        \registers[16][28] ), .B2(n1950), .ZN(n1055) );
  OAI221_X1 U1097 ( .B1(n1959), .B2(n2459), .C1(n1956), .C2(n2427), .A(n1072), 
        .ZN(n1071) );
  AOI22_X1 U1098 ( .A1(\registers[17][29] ), .A2(n1953), .B1(
        \registers[16][29] ), .B2(n1950), .ZN(n1072) );
  OAI221_X1 U1099 ( .B1(n1959), .B2(n2458), .C1(n1956), .C2(n2426), .A(n1089), 
        .ZN(n1088) );
  AOI22_X1 U1100 ( .A1(\registers[17][30] ), .A2(n1953), .B1(
        \registers[16][30] ), .B2(n1950), .ZN(n1089) );
  OAI221_X1 U1101 ( .B1(n1959), .B2(n2457), .C1(n1956), .C2(n2425), .A(n1106), 
        .ZN(n1105) );
  AOI22_X1 U1102 ( .A1(\registers[17][31] ), .A2(n1953), .B1(
        \registers[16][31] ), .B2(n1950), .ZN(n1106) );
  OAI221_X1 U1103 ( .B1(n1904), .B2(n2200), .C1(n1901), .C2(n2264), .A(n575), 
        .ZN(n569) );
  AOI22_X1 U1104 ( .A1(\registers[3][0] ), .A2(n1898), .B1(\registers[6][0] ), 
        .B2(n1895), .ZN(n575) );
  OAI221_X1 U1105 ( .B1(n1904), .B2(n2199), .C1(n1901), .C2(n2263), .A(n602), 
        .ZN(n600) );
  AOI22_X1 U1106 ( .A1(\registers[3][1] ), .A2(n1898), .B1(\registers[6][1] ), 
        .B2(n1895), .ZN(n602) );
  OAI221_X1 U1107 ( .B1(n1904), .B2(n2198), .C1(n1901), .C2(n2262), .A(n619), 
        .ZN(n617) );
  AOI22_X1 U1108 ( .A1(\registers[3][2] ), .A2(n1898), .B1(\registers[6][2] ), 
        .B2(n1895), .ZN(n619) );
  OAI221_X1 U1109 ( .B1(n1904), .B2(n2197), .C1(n1901), .C2(n2261), .A(n636), 
        .ZN(n634) );
  AOI22_X1 U1110 ( .A1(\registers[3][3] ), .A2(n1898), .B1(\registers[6][3] ), 
        .B2(n1895), .ZN(n636) );
  OAI221_X1 U1111 ( .B1(n1904), .B2(n2196), .C1(n1901), .C2(n2260), .A(n653), 
        .ZN(n651) );
  AOI22_X1 U1112 ( .A1(\registers[3][4] ), .A2(n1898), .B1(\registers[6][4] ), 
        .B2(n1895), .ZN(n653) );
  OAI221_X1 U1113 ( .B1(n1904), .B2(n2195), .C1(n1901), .C2(n2259), .A(n670), 
        .ZN(n668) );
  AOI22_X1 U1114 ( .A1(\registers[3][5] ), .A2(n1898), .B1(\registers[6][5] ), 
        .B2(n1895), .ZN(n670) );
  OAI221_X1 U1115 ( .B1(n1904), .B2(n2194), .C1(n1901), .C2(n2258), .A(n687), 
        .ZN(n685) );
  AOI22_X1 U1116 ( .A1(\registers[3][6] ), .A2(n1898), .B1(\registers[6][6] ), 
        .B2(n1895), .ZN(n687) );
  OAI221_X1 U1117 ( .B1(n1904), .B2(n2193), .C1(n1901), .C2(n2257), .A(n704), 
        .ZN(n702) );
  AOI22_X1 U1118 ( .A1(\registers[3][7] ), .A2(n1898), .B1(\registers[6][7] ), 
        .B2(n1895), .ZN(n704) );
  OAI221_X1 U1119 ( .B1(n2200), .B2(n1811), .C1(n2264), .C2(n1808), .A(n1162), 
        .ZN(n1156) );
  AOI22_X1 U1120 ( .A1(n1805), .A2(\registers[3][0] ), .B1(n1800), .B2(
        \registers[6][0] ), .ZN(n1162) );
  OAI221_X1 U1121 ( .B1(n2199), .B2(n1811), .C1(n2263), .C2(n1808), .A(n1189), 
        .ZN(n1187) );
  AOI22_X1 U1122 ( .A1(n1805), .A2(\registers[3][1] ), .B1(n1800), .B2(
        \registers[6][1] ), .ZN(n1189) );
  OAI221_X1 U1123 ( .B1(n2198), .B2(n1811), .C1(n2262), .C2(n1808), .A(n1206), 
        .ZN(n1204) );
  AOI22_X1 U1124 ( .A1(n1805), .A2(\registers[3][2] ), .B1(n1800), .B2(
        \registers[6][2] ), .ZN(n1206) );
  OAI221_X1 U1125 ( .B1(n2197), .B2(n1811), .C1(n2261), .C2(n1808), .A(n1223), 
        .ZN(n1221) );
  AOI22_X1 U1126 ( .A1(n1805), .A2(\registers[3][3] ), .B1(n1800), .B2(
        \registers[6][3] ), .ZN(n1223) );
  OAI221_X1 U1127 ( .B1(n2196), .B2(n1811), .C1(n2260), .C2(n1808), .A(n1240), 
        .ZN(n1238) );
  AOI22_X1 U1128 ( .A1(n1805), .A2(\registers[3][4] ), .B1(n1800), .B2(
        \registers[6][4] ), .ZN(n1240) );
  OAI221_X1 U1129 ( .B1(n2195), .B2(n1811), .C1(n2259), .C2(n1808), .A(n1257), 
        .ZN(n1255) );
  AOI22_X1 U1130 ( .A1(n1805), .A2(\registers[3][5] ), .B1(n1800), .B2(
        \registers[6][5] ), .ZN(n1257) );
  OAI221_X1 U1131 ( .B1(n2194), .B2(n1811), .C1(n2258), .C2(n1808), .A(n1274), 
        .ZN(n1272) );
  AOI22_X1 U1132 ( .A1(n1805), .A2(\registers[3][6] ), .B1(n1800), .B2(
        \registers[6][6] ), .ZN(n1274) );
  OAI221_X1 U1133 ( .B1(n2193), .B2(n1811), .C1(n2257), .C2(n1808), .A(n1291), 
        .ZN(n1289) );
  AOI22_X1 U1134 ( .A1(n1805), .A2(\registers[3][7] ), .B1(n1800), .B2(
        \registers[6][7] ), .ZN(n1291) );
  OAI221_X1 U1135 ( .B1(n2192), .B2(n1810), .C1(n2256), .C2(n1807), .A(n1308), 
        .ZN(n1306) );
  AOI22_X1 U1136 ( .A1(n1804), .A2(\registers[3][8] ), .B1(n1800), .B2(
        \registers[6][8] ), .ZN(n1308) );
  OAI221_X1 U1137 ( .B1(n2191), .B2(n1810), .C1(n2255), .C2(n1807), .A(n1325), 
        .ZN(n1323) );
  AOI22_X1 U1138 ( .A1(n1804), .A2(\registers[3][9] ), .B1(n1800), .B2(
        \registers[6][9] ), .ZN(n1325) );
  OAI221_X1 U1139 ( .B1(n2190), .B2(n1810), .C1(n2254), .C2(n1807), .A(n1342), 
        .ZN(n1340) );
  AOI22_X1 U1140 ( .A1(n1804), .A2(\registers[3][10] ), .B1(n1800), .B2(
        \registers[6][10] ), .ZN(n1342) );
  OAI221_X1 U1141 ( .B1(n2189), .B2(n1810), .C1(n2253), .C2(n1807), .A(n1359), 
        .ZN(n1357) );
  AOI22_X1 U1142 ( .A1(n1804), .A2(\registers[3][11] ), .B1(n1800), .B2(
        \registers[6][11] ), .ZN(n1359) );
  OAI221_X1 U1143 ( .B1(n2188), .B2(n1810), .C1(n2252), .C2(n1807), .A(n1376), 
        .ZN(n1374) );
  AOI22_X1 U1144 ( .A1(n1804), .A2(\registers[3][12] ), .B1(n1801), .B2(
        \registers[6][12] ), .ZN(n1376) );
  OAI221_X1 U1145 ( .B1(n2187), .B2(n1810), .C1(n2251), .C2(n1807), .A(n1393), 
        .ZN(n1391) );
  AOI22_X1 U1146 ( .A1(n1804), .A2(\registers[3][13] ), .B1(n1801), .B2(
        \registers[6][13] ), .ZN(n1393) );
  OAI221_X1 U1147 ( .B1(n2186), .B2(n1810), .C1(n2250), .C2(n1807), .A(n1410), 
        .ZN(n1408) );
  AOI22_X1 U1148 ( .A1(n1804), .A2(\registers[3][14] ), .B1(n1801), .B2(
        \registers[6][14] ), .ZN(n1410) );
  OAI221_X1 U1149 ( .B1(n2185), .B2(n1810), .C1(n2249), .C2(n1807), .A(n1427), 
        .ZN(n1425) );
  AOI22_X1 U1150 ( .A1(n1804), .A2(\registers[3][15] ), .B1(n1801), .B2(
        \registers[6][15] ), .ZN(n1427) );
  OAI221_X1 U1151 ( .B1(n2184), .B2(n1810), .C1(n2248), .C2(n1807), .A(n1444), 
        .ZN(n1442) );
  AOI22_X1 U1152 ( .A1(n1804), .A2(\registers[3][16] ), .B1(n1801), .B2(
        \registers[6][16] ), .ZN(n1444) );
  OAI221_X1 U1153 ( .B1(n2183), .B2(n1810), .C1(n2247), .C2(n1807), .A(n1461), 
        .ZN(n1459) );
  AOI22_X1 U1154 ( .A1(n1804), .A2(\registers[3][17] ), .B1(n1801), .B2(
        \registers[6][17] ), .ZN(n1461) );
  OAI221_X1 U1155 ( .B1(n2182), .B2(n1810), .C1(n2246), .C2(n1807), .A(n1478), 
        .ZN(n1476) );
  AOI22_X1 U1156 ( .A1(n1804), .A2(\registers[3][18] ), .B1(n1801), .B2(
        \registers[6][18] ), .ZN(n1478) );
  OAI221_X1 U1157 ( .B1(n2181), .B2(n1810), .C1(n2245), .C2(n1807), .A(n1495), 
        .ZN(n1493) );
  AOI22_X1 U1158 ( .A1(n1804), .A2(\registers[3][19] ), .B1(n1801), .B2(
        \registers[6][19] ), .ZN(n1495) );
  OAI221_X1 U1159 ( .B1(n2180), .B2(n1809), .C1(n2244), .C2(n1806), .A(n1512), 
        .ZN(n1510) );
  AOI22_X1 U1160 ( .A1(n1803), .A2(\registers[3][20] ), .B1(n1801), .B2(
        \registers[6][20] ), .ZN(n1512) );
  OAI221_X1 U1161 ( .B1(n2179), .B2(n1809), .C1(n2243), .C2(n1806), .A(n1529), 
        .ZN(n1527) );
  AOI22_X1 U1162 ( .A1(n1803), .A2(\registers[3][21] ), .B1(n1801), .B2(
        \registers[6][21] ), .ZN(n1529) );
  OAI221_X1 U1163 ( .B1(n2178), .B2(n1809), .C1(n2242), .C2(n1806), .A(n1546), 
        .ZN(n1544) );
  AOI22_X1 U1164 ( .A1(n1803), .A2(\registers[3][22] ), .B1(n1801), .B2(
        \registers[6][22] ), .ZN(n1546) );
  OAI221_X1 U1165 ( .B1(n2177), .B2(n1809), .C1(n2241), .C2(n1806), .A(n1563), 
        .ZN(n1561) );
  AOI22_X1 U1166 ( .A1(n1803), .A2(\registers[3][23] ), .B1(n1801), .B2(
        \registers[6][23] ), .ZN(n1563) );
  OAI221_X1 U1167 ( .B1(n2176), .B2(n1809), .C1(n2240), .C2(n1806), .A(n1580), 
        .ZN(n1578) );
  AOI22_X1 U1168 ( .A1(n1803), .A2(\registers[3][24] ), .B1(n1802), .B2(
        \registers[6][24] ), .ZN(n1580) );
  OAI221_X1 U1169 ( .B1(n2175), .B2(n1809), .C1(n2239), .C2(n1806), .A(n1597), 
        .ZN(n1595) );
  AOI22_X1 U1170 ( .A1(n1803), .A2(\registers[3][25] ), .B1(n1802), .B2(
        \registers[6][25] ), .ZN(n1597) );
  OAI221_X1 U1171 ( .B1(n2174), .B2(n1809), .C1(n2238), .C2(n1806), .A(n1614), 
        .ZN(n1612) );
  AOI22_X1 U1172 ( .A1(n1803), .A2(\registers[3][26] ), .B1(n1802), .B2(
        \registers[6][26] ), .ZN(n1614) );
  OAI221_X1 U1173 ( .B1(n2173), .B2(n1809), .C1(n2237), .C2(n1806), .A(n1631), 
        .ZN(n1629) );
  AOI22_X1 U1174 ( .A1(n1803), .A2(\registers[3][27] ), .B1(n1802), .B2(
        \registers[6][27] ), .ZN(n1631) );
  OAI221_X1 U1175 ( .B1(n2172), .B2(n1809), .C1(n2236), .C2(n1806), .A(n1648), 
        .ZN(n1646) );
  AOI22_X1 U1176 ( .A1(n1803), .A2(\registers[3][28] ), .B1(n1802), .B2(
        \registers[6][28] ), .ZN(n1648) );
  OAI221_X1 U1177 ( .B1(n2171), .B2(n1809), .C1(n2235), .C2(n1806), .A(n1665), 
        .ZN(n1663) );
  AOI22_X1 U1178 ( .A1(n1803), .A2(\registers[3][29] ), .B1(n1802), .B2(
        \registers[6][29] ), .ZN(n1665) );
  OAI221_X1 U1179 ( .B1(n2170), .B2(n1809), .C1(n2234), .C2(n1806), .A(n1682), 
        .ZN(n1680) );
  AOI22_X1 U1180 ( .A1(n1803), .A2(\registers[3][30] ), .B1(n1802), .B2(
        \registers[6][30] ), .ZN(n1682) );
  OAI221_X1 U1181 ( .B1(n2169), .B2(n1809), .C1(n2233), .C2(n1806), .A(n1709), 
        .ZN(n1705) );
  AOI22_X1 U1182 ( .A1(n1803), .A2(\registers[3][31] ), .B1(n1802), .B2(
        \registers[6][31] ), .ZN(n1709) );
  OAI221_X1 U1183 ( .B1(n1903), .B2(n2192), .C1(n1900), .C2(n2256), .A(n721), 
        .ZN(n719) );
  AOI22_X1 U1184 ( .A1(\registers[3][8] ), .A2(n1897), .B1(\registers[6][8] ), 
        .B2(n1894), .ZN(n721) );
  OAI221_X1 U1185 ( .B1(n1903), .B2(n2191), .C1(n1900), .C2(n2255), .A(n738), 
        .ZN(n736) );
  AOI22_X1 U1186 ( .A1(\registers[3][9] ), .A2(n1897), .B1(\registers[6][9] ), 
        .B2(n1894), .ZN(n738) );
  OAI221_X1 U1187 ( .B1(n1903), .B2(n2190), .C1(n1900), .C2(n2254), .A(n755), 
        .ZN(n753) );
  AOI22_X1 U1188 ( .A1(\registers[3][10] ), .A2(n1897), .B1(\registers[6][10] ), .B2(n1894), .ZN(n755) );
  OAI221_X1 U1189 ( .B1(n1903), .B2(n2189), .C1(n1900), .C2(n2253), .A(n772), 
        .ZN(n770) );
  AOI22_X1 U1190 ( .A1(\registers[3][11] ), .A2(n1897), .B1(\registers[6][11] ), .B2(n1894), .ZN(n772) );
  OAI221_X1 U1191 ( .B1(n1903), .B2(n2188), .C1(n1900), .C2(n2252), .A(n789), 
        .ZN(n787) );
  AOI22_X1 U1192 ( .A1(\registers[3][12] ), .A2(n1897), .B1(\registers[6][12] ), .B2(n1894), .ZN(n789) );
  OAI221_X1 U1193 ( .B1(n1903), .B2(n2187), .C1(n1900), .C2(n2251), .A(n806), 
        .ZN(n804) );
  AOI22_X1 U1194 ( .A1(\registers[3][13] ), .A2(n1897), .B1(\registers[6][13] ), .B2(n1894), .ZN(n806) );
  OAI221_X1 U1195 ( .B1(n1903), .B2(n2186), .C1(n1900), .C2(n2250), .A(n823), 
        .ZN(n821) );
  AOI22_X1 U1196 ( .A1(\registers[3][14] ), .A2(n1897), .B1(\registers[6][14] ), .B2(n1894), .ZN(n823) );
  OAI221_X1 U1197 ( .B1(n1903), .B2(n2185), .C1(n1900), .C2(n2249), .A(n840), 
        .ZN(n838) );
  AOI22_X1 U1198 ( .A1(\registers[3][15] ), .A2(n1897), .B1(\registers[6][15] ), .B2(n1894), .ZN(n840) );
  OAI221_X1 U1199 ( .B1(n1903), .B2(n2184), .C1(n1900), .C2(n2248), .A(n857), 
        .ZN(n855) );
  AOI22_X1 U1200 ( .A1(\registers[3][16] ), .A2(n1897), .B1(\registers[6][16] ), .B2(n1894), .ZN(n857) );
  OAI221_X1 U1201 ( .B1(n1903), .B2(n2183), .C1(n1900), .C2(n2247), .A(n874), 
        .ZN(n872) );
  AOI22_X1 U1202 ( .A1(\registers[3][17] ), .A2(n1897), .B1(\registers[6][17] ), .B2(n1894), .ZN(n874) );
  OAI221_X1 U1203 ( .B1(n1903), .B2(n2182), .C1(n1900), .C2(n2246), .A(n891), 
        .ZN(n889) );
  AOI22_X1 U1204 ( .A1(\registers[3][18] ), .A2(n1897), .B1(\registers[6][18] ), .B2(n1894), .ZN(n891) );
  OAI221_X1 U1205 ( .B1(n1903), .B2(n2181), .C1(n1900), .C2(n2245), .A(n908), 
        .ZN(n906) );
  AOI22_X1 U1206 ( .A1(\registers[3][19] ), .A2(n1897), .B1(\registers[6][19] ), .B2(n1894), .ZN(n908) );
  OAI221_X1 U1207 ( .B1(n1902), .B2(n2180), .C1(n1899), .C2(n2244), .A(n925), 
        .ZN(n923) );
  AOI22_X1 U1208 ( .A1(\registers[3][20] ), .A2(n1896), .B1(\registers[6][20] ), .B2(n1893), .ZN(n925) );
  OAI221_X1 U1209 ( .B1(n1902), .B2(n2179), .C1(n1899), .C2(n2243), .A(n942), 
        .ZN(n940) );
  AOI22_X1 U1210 ( .A1(\registers[3][21] ), .A2(n1896), .B1(\registers[6][21] ), .B2(n1893), .ZN(n942) );
  OAI221_X1 U1211 ( .B1(n1902), .B2(n2178), .C1(n1899), .C2(n2242), .A(n959), 
        .ZN(n957) );
  AOI22_X1 U1212 ( .A1(\registers[3][22] ), .A2(n1896), .B1(\registers[6][22] ), .B2(n1893), .ZN(n959) );
  OAI221_X1 U1213 ( .B1(n1902), .B2(n2177), .C1(n1899), .C2(n2241), .A(n976), 
        .ZN(n974) );
  AOI22_X1 U1214 ( .A1(\registers[3][23] ), .A2(n1896), .B1(\registers[6][23] ), .B2(n1893), .ZN(n976) );
  OAI221_X1 U1215 ( .B1(n1902), .B2(n2176), .C1(n1899), .C2(n2240), .A(n993), 
        .ZN(n991) );
  AOI22_X1 U1216 ( .A1(\registers[3][24] ), .A2(n1896), .B1(\registers[6][24] ), .B2(n1893), .ZN(n993) );
  OAI221_X1 U1217 ( .B1(n1902), .B2(n2175), .C1(n1899), .C2(n2239), .A(n1010), 
        .ZN(n1008) );
  AOI22_X1 U1218 ( .A1(\registers[3][25] ), .A2(n1896), .B1(\registers[6][25] ), .B2(n1893), .ZN(n1010) );
  OAI221_X1 U1219 ( .B1(n1902), .B2(n2174), .C1(n1899), .C2(n2238), .A(n1027), 
        .ZN(n1025) );
  AOI22_X1 U1220 ( .A1(\registers[3][26] ), .A2(n1896), .B1(\registers[6][26] ), .B2(n1893), .ZN(n1027) );
  OAI221_X1 U1221 ( .B1(n1902), .B2(n2173), .C1(n1899), .C2(n2237), .A(n1044), 
        .ZN(n1042) );
  AOI22_X1 U1222 ( .A1(\registers[3][27] ), .A2(n1896), .B1(\registers[6][27] ), .B2(n1893), .ZN(n1044) );
  OAI221_X1 U1223 ( .B1(n1902), .B2(n2172), .C1(n1899), .C2(n2236), .A(n1061), 
        .ZN(n1059) );
  AOI22_X1 U1224 ( .A1(\registers[3][28] ), .A2(n1896), .B1(\registers[6][28] ), .B2(n1893), .ZN(n1061) );
  OAI221_X1 U1225 ( .B1(n1902), .B2(n2171), .C1(n1899), .C2(n2235), .A(n1078), 
        .ZN(n1076) );
  AOI22_X1 U1226 ( .A1(\registers[3][29] ), .A2(n1896), .B1(\registers[6][29] ), .B2(n1893), .ZN(n1078) );
  OAI221_X1 U1227 ( .B1(n1902), .B2(n2170), .C1(n1899), .C2(n2234), .A(n1095), 
        .ZN(n1093) );
  AOI22_X1 U1228 ( .A1(\registers[3][30] ), .A2(n1896), .B1(\registers[6][30] ), .B2(n1893), .ZN(n1095) );
  OAI221_X1 U1229 ( .B1(n1902), .B2(n2169), .C1(n1899), .C2(n2233), .A(n1122), 
        .ZN(n1118) );
  AOI22_X1 U1230 ( .A1(\registers[3][31] ), .A2(n1896), .B1(\registers[6][31] ), .B2(n1893), .ZN(n1122) );
  AOI22_X1 U1231 ( .A1(\registers[23][0] ), .A2(n1943), .B1(\registers[22][0] ), .B2(n1940), .ZN(n555) );
  AOI22_X1 U1232 ( .A1(\registers[25][0] ), .A2(n1931), .B1(\registers[24][0] ), .B2(n1928), .ZN(n560) );
  AOI22_X1 U1233 ( .A1(\registers[31][0] ), .A2(n1919), .B1(\registers[30][0] ), .B2(n1916), .ZN(n565) );
  AOI22_X1 U1234 ( .A1(\registers[23][1] ), .A2(n1943), .B1(\registers[22][1] ), .B2(n1940), .ZN(n597) );
  AOI22_X1 U1235 ( .A1(\registers[25][1] ), .A2(n1931), .B1(\registers[24][1] ), .B2(n1928), .ZN(n598) );
  AOI22_X1 U1236 ( .A1(\registers[31][1] ), .A2(n1919), .B1(\registers[30][1] ), .B2(n1916), .ZN(n599) );
  AOI22_X1 U1237 ( .A1(\registers[23][2] ), .A2(n1943), .B1(\registers[22][2] ), .B2(n1940), .ZN(n614) );
  AOI22_X1 U1238 ( .A1(\registers[25][2] ), .A2(n1931), .B1(\registers[24][2] ), .B2(n1928), .ZN(n615) );
  AOI22_X1 U1239 ( .A1(\registers[31][2] ), .A2(n1919), .B1(\registers[30][2] ), .B2(n1916), .ZN(n616) );
  AOI22_X1 U1240 ( .A1(\registers[23][3] ), .A2(n1943), .B1(\registers[22][3] ), .B2(n1940), .ZN(n631) );
  AOI22_X1 U1241 ( .A1(\registers[25][3] ), .A2(n1931), .B1(\registers[24][3] ), .B2(n1928), .ZN(n632) );
  AOI22_X1 U1242 ( .A1(\registers[31][3] ), .A2(n1919), .B1(\registers[30][3] ), .B2(n1916), .ZN(n633) );
  AOI22_X1 U1243 ( .A1(\registers[23][4] ), .A2(n1943), .B1(\registers[22][4] ), .B2(n1940), .ZN(n648) );
  AOI22_X1 U1244 ( .A1(\registers[25][4] ), .A2(n1931), .B1(\registers[24][4] ), .B2(n1928), .ZN(n649) );
  AOI22_X1 U1245 ( .A1(\registers[31][4] ), .A2(n1919), .B1(\registers[30][4] ), .B2(n1916), .ZN(n650) );
  AOI22_X1 U1246 ( .A1(\registers[23][5] ), .A2(n1943), .B1(\registers[22][5] ), .B2(n1940), .ZN(n665) );
  AOI22_X1 U1247 ( .A1(\registers[25][5] ), .A2(n1931), .B1(\registers[24][5] ), .B2(n1928), .ZN(n666) );
  AOI22_X1 U1248 ( .A1(\registers[31][5] ), .A2(n1919), .B1(\registers[30][5] ), .B2(n1916), .ZN(n667) );
  AOI22_X1 U1249 ( .A1(\registers[23][6] ), .A2(n1943), .B1(\registers[22][6] ), .B2(n1940), .ZN(n682) );
  AOI22_X1 U1250 ( .A1(\registers[25][6] ), .A2(n1931), .B1(\registers[24][6] ), .B2(n1928), .ZN(n683) );
  AOI22_X1 U1251 ( .A1(\registers[31][6] ), .A2(n1919), .B1(\registers[30][6] ), .B2(n1916), .ZN(n684) );
  AOI22_X1 U1252 ( .A1(\registers[23][7] ), .A2(n1943), .B1(\registers[22][7] ), .B2(n1940), .ZN(n699) );
  AOI22_X1 U1253 ( .A1(\registers[25][7] ), .A2(n1931), .B1(\registers[24][7] ), .B2(n1928), .ZN(n700) );
  AOI22_X1 U1254 ( .A1(\registers[31][7] ), .A2(n1919), .B1(\registers[30][7] ), .B2(n1916), .ZN(n701) );
  AOI22_X1 U1255 ( .A1(n1850), .A2(\registers[23][0] ), .B1(n1845), .B2(
        \registers[22][0] ), .ZN(n1142) );
  AOI22_X1 U1256 ( .A1(n1838), .A2(\registers[25][0] ), .B1(n1833), .B2(
        \registers[24][0] ), .ZN(n1147) );
  AOI22_X1 U1257 ( .A1(n1826), .A2(\registers[31][0] ), .B1(n1821), .B2(
        \registers[30][0] ), .ZN(n1152) );
  AOI22_X1 U1258 ( .A1(n1850), .A2(\registers[23][1] ), .B1(n1845), .B2(
        \registers[22][1] ), .ZN(n1184) );
  AOI22_X1 U1259 ( .A1(n1838), .A2(\registers[25][1] ), .B1(n1833), .B2(
        \registers[24][1] ), .ZN(n1185) );
  AOI22_X1 U1260 ( .A1(n1826), .A2(\registers[31][1] ), .B1(n1821), .B2(
        \registers[30][1] ), .ZN(n1186) );
  AOI22_X1 U1261 ( .A1(n1850), .A2(\registers[23][2] ), .B1(n1845), .B2(
        \registers[22][2] ), .ZN(n1201) );
  AOI22_X1 U1262 ( .A1(n1838), .A2(\registers[25][2] ), .B1(n1833), .B2(
        \registers[24][2] ), .ZN(n1202) );
  AOI22_X1 U1263 ( .A1(n1826), .A2(\registers[31][2] ), .B1(n1821), .B2(
        \registers[30][2] ), .ZN(n1203) );
  AOI22_X1 U1264 ( .A1(n1850), .A2(\registers[23][3] ), .B1(n1845), .B2(
        \registers[22][3] ), .ZN(n1218) );
  AOI22_X1 U1265 ( .A1(n1838), .A2(\registers[25][3] ), .B1(n1833), .B2(
        \registers[24][3] ), .ZN(n1219) );
  AOI22_X1 U1266 ( .A1(n1826), .A2(\registers[31][3] ), .B1(n1821), .B2(
        \registers[30][3] ), .ZN(n1220) );
  AOI22_X1 U1267 ( .A1(n1850), .A2(\registers[23][4] ), .B1(n1845), .B2(
        \registers[22][4] ), .ZN(n1235) );
  AOI22_X1 U1268 ( .A1(n1838), .A2(\registers[25][4] ), .B1(n1833), .B2(
        \registers[24][4] ), .ZN(n1236) );
  AOI22_X1 U1269 ( .A1(n1826), .A2(\registers[31][4] ), .B1(n1821), .B2(
        \registers[30][4] ), .ZN(n1237) );
  AOI22_X1 U1270 ( .A1(n1850), .A2(\registers[23][5] ), .B1(n1845), .B2(
        \registers[22][5] ), .ZN(n1252) );
  AOI22_X1 U1271 ( .A1(n1838), .A2(\registers[25][5] ), .B1(n1833), .B2(
        \registers[24][5] ), .ZN(n1253) );
  AOI22_X1 U1272 ( .A1(n1826), .A2(\registers[31][5] ), .B1(n1821), .B2(
        \registers[30][5] ), .ZN(n1254) );
  AOI22_X1 U1273 ( .A1(n1850), .A2(\registers[23][6] ), .B1(n1845), .B2(
        \registers[22][6] ), .ZN(n1269) );
  AOI22_X1 U1274 ( .A1(n1838), .A2(\registers[25][6] ), .B1(n1833), .B2(
        \registers[24][6] ), .ZN(n1270) );
  AOI22_X1 U1275 ( .A1(n1826), .A2(\registers[31][6] ), .B1(n1821), .B2(
        \registers[30][6] ), .ZN(n1271) );
  AOI22_X1 U1276 ( .A1(n1850), .A2(\registers[23][7] ), .B1(n1845), .B2(
        \registers[22][7] ), .ZN(n1286) );
  AOI22_X1 U1277 ( .A1(n1838), .A2(\registers[25][7] ), .B1(n1833), .B2(
        \registers[24][7] ), .ZN(n1287) );
  AOI22_X1 U1278 ( .A1(n1826), .A2(\registers[31][7] ), .B1(n1821), .B2(
        \registers[30][7] ), .ZN(n1288) );
  AOI22_X1 U1279 ( .A1(n1849), .A2(\registers[23][8] ), .B1(n1845), .B2(
        \registers[22][8] ), .ZN(n1303) );
  AOI22_X1 U1280 ( .A1(n1837), .A2(\registers[25][8] ), .B1(n1833), .B2(
        \registers[24][8] ), .ZN(n1304) );
  AOI22_X1 U1281 ( .A1(n1825), .A2(\registers[31][8] ), .B1(n1821), .B2(
        \registers[30][8] ), .ZN(n1305) );
  AOI22_X1 U1282 ( .A1(n1849), .A2(\registers[23][9] ), .B1(n1845), .B2(
        \registers[22][9] ), .ZN(n1320) );
  AOI22_X1 U1283 ( .A1(n1837), .A2(\registers[25][9] ), .B1(n1833), .B2(
        \registers[24][9] ), .ZN(n1321) );
  AOI22_X1 U1284 ( .A1(n1825), .A2(\registers[31][9] ), .B1(n1821), .B2(
        \registers[30][9] ), .ZN(n1322) );
  AOI22_X1 U1285 ( .A1(n1849), .A2(\registers[23][10] ), .B1(n1845), .B2(
        \registers[22][10] ), .ZN(n1337) );
  AOI22_X1 U1286 ( .A1(n1837), .A2(\registers[25][10] ), .B1(n1833), .B2(
        \registers[24][10] ), .ZN(n1338) );
  AOI22_X1 U1287 ( .A1(n1825), .A2(\registers[31][10] ), .B1(n1821), .B2(
        \registers[30][10] ), .ZN(n1339) );
  AOI22_X1 U1288 ( .A1(n1849), .A2(\registers[23][11] ), .B1(n1845), .B2(
        \registers[22][11] ), .ZN(n1354) );
  AOI22_X1 U1289 ( .A1(n1837), .A2(\registers[25][11] ), .B1(n1833), .B2(
        \registers[24][11] ), .ZN(n1355) );
  AOI22_X1 U1290 ( .A1(n1825), .A2(\registers[31][11] ), .B1(n1821), .B2(
        \registers[30][11] ), .ZN(n1356) );
  AOI22_X1 U1291 ( .A1(n1849), .A2(\registers[23][12] ), .B1(n1846), .B2(
        \registers[22][12] ), .ZN(n1371) );
  AOI22_X1 U1292 ( .A1(n1837), .A2(\registers[25][12] ), .B1(n1834), .B2(
        \registers[24][12] ), .ZN(n1372) );
  AOI22_X1 U1293 ( .A1(n1825), .A2(\registers[31][12] ), .B1(n1822), .B2(
        \registers[30][12] ), .ZN(n1373) );
  AOI22_X1 U1294 ( .A1(n1849), .A2(\registers[23][13] ), .B1(n1846), .B2(
        \registers[22][13] ), .ZN(n1388) );
  AOI22_X1 U1295 ( .A1(n1837), .A2(\registers[25][13] ), .B1(n1834), .B2(
        \registers[24][13] ), .ZN(n1389) );
  AOI22_X1 U1296 ( .A1(n1825), .A2(\registers[31][13] ), .B1(n1822), .B2(
        \registers[30][13] ), .ZN(n1390) );
  AOI22_X1 U1297 ( .A1(n1849), .A2(\registers[23][14] ), .B1(n1846), .B2(
        \registers[22][14] ), .ZN(n1405) );
  AOI22_X1 U1298 ( .A1(n1837), .A2(\registers[25][14] ), .B1(n1834), .B2(
        \registers[24][14] ), .ZN(n1406) );
  AOI22_X1 U1299 ( .A1(n1825), .A2(\registers[31][14] ), .B1(n1822), .B2(
        \registers[30][14] ), .ZN(n1407) );
  AOI22_X1 U1300 ( .A1(n1849), .A2(\registers[23][15] ), .B1(n1846), .B2(
        \registers[22][15] ), .ZN(n1422) );
  AOI22_X1 U1301 ( .A1(n1837), .A2(\registers[25][15] ), .B1(n1834), .B2(
        \registers[24][15] ), .ZN(n1423) );
  AOI22_X1 U1302 ( .A1(n1825), .A2(\registers[31][15] ), .B1(n1822), .B2(
        \registers[30][15] ), .ZN(n1424) );
  AOI22_X1 U1303 ( .A1(n1849), .A2(\registers[23][16] ), .B1(n1846), .B2(
        \registers[22][16] ), .ZN(n1439) );
  AOI22_X1 U1304 ( .A1(n1837), .A2(\registers[25][16] ), .B1(n1834), .B2(
        \registers[24][16] ), .ZN(n1440) );
  AOI22_X1 U1305 ( .A1(n1825), .A2(\registers[31][16] ), .B1(n1822), .B2(
        \registers[30][16] ), .ZN(n1441) );
  AOI22_X1 U1306 ( .A1(n1849), .A2(\registers[23][17] ), .B1(n1846), .B2(
        \registers[22][17] ), .ZN(n1456) );
  AOI22_X1 U1307 ( .A1(n1837), .A2(\registers[25][17] ), .B1(n1834), .B2(
        \registers[24][17] ), .ZN(n1457) );
  AOI22_X1 U1308 ( .A1(n1825), .A2(\registers[31][17] ), .B1(n1822), .B2(
        \registers[30][17] ), .ZN(n1458) );
  AOI22_X1 U1309 ( .A1(n1849), .A2(\registers[23][18] ), .B1(n1846), .B2(
        \registers[22][18] ), .ZN(n1473) );
  AOI22_X1 U1310 ( .A1(n1837), .A2(\registers[25][18] ), .B1(n1834), .B2(
        \registers[24][18] ), .ZN(n1474) );
  AOI22_X1 U1311 ( .A1(n1825), .A2(\registers[31][18] ), .B1(n1822), .B2(
        \registers[30][18] ), .ZN(n1475) );
  AOI22_X1 U1312 ( .A1(n1849), .A2(\registers[23][19] ), .B1(n1846), .B2(
        \registers[22][19] ), .ZN(n1490) );
  AOI22_X1 U1313 ( .A1(n1837), .A2(\registers[25][19] ), .B1(n1834), .B2(
        \registers[24][19] ), .ZN(n1491) );
  AOI22_X1 U1314 ( .A1(n1825), .A2(\registers[31][19] ), .B1(n1822), .B2(
        \registers[30][19] ), .ZN(n1492) );
  AOI22_X1 U1315 ( .A1(n1848), .A2(\registers[23][20] ), .B1(n1846), .B2(
        \registers[22][20] ), .ZN(n1507) );
  AOI22_X1 U1316 ( .A1(n1836), .A2(\registers[25][20] ), .B1(n1834), .B2(
        \registers[24][20] ), .ZN(n1508) );
  AOI22_X1 U1317 ( .A1(n1824), .A2(\registers[31][20] ), .B1(n1822), .B2(
        \registers[30][20] ), .ZN(n1509) );
  AOI22_X1 U1318 ( .A1(n1848), .A2(\registers[23][21] ), .B1(n1846), .B2(
        \registers[22][21] ), .ZN(n1524) );
  AOI22_X1 U1319 ( .A1(n1836), .A2(\registers[25][21] ), .B1(n1834), .B2(
        \registers[24][21] ), .ZN(n1525) );
  AOI22_X1 U1320 ( .A1(n1824), .A2(\registers[31][21] ), .B1(n1822), .B2(
        \registers[30][21] ), .ZN(n1526) );
  AOI22_X1 U1321 ( .A1(n1848), .A2(\registers[23][22] ), .B1(n1846), .B2(
        \registers[22][22] ), .ZN(n1541) );
  AOI22_X1 U1322 ( .A1(n1836), .A2(\registers[25][22] ), .B1(n1834), .B2(
        \registers[24][22] ), .ZN(n1542) );
  AOI22_X1 U1323 ( .A1(n1824), .A2(\registers[31][22] ), .B1(n1822), .B2(
        \registers[30][22] ), .ZN(n1543) );
  AOI22_X1 U1324 ( .A1(n1848), .A2(\registers[23][23] ), .B1(n1846), .B2(
        \registers[22][23] ), .ZN(n1558) );
  AOI22_X1 U1325 ( .A1(n1836), .A2(\registers[25][23] ), .B1(n1834), .B2(
        \registers[24][23] ), .ZN(n1559) );
  AOI22_X1 U1326 ( .A1(n1824), .A2(\registers[31][23] ), .B1(n1822), .B2(
        \registers[30][23] ), .ZN(n1560) );
  AOI22_X1 U1327 ( .A1(n1848), .A2(\registers[23][24] ), .B1(n1847), .B2(
        \registers[22][24] ), .ZN(n1575) );
  AOI22_X1 U1328 ( .A1(n1836), .A2(\registers[25][24] ), .B1(n1835), .B2(
        \registers[24][24] ), .ZN(n1576) );
  AOI22_X1 U1329 ( .A1(n1824), .A2(\registers[31][24] ), .B1(n1823), .B2(
        \registers[30][24] ), .ZN(n1577) );
  AOI22_X1 U1330 ( .A1(n1848), .A2(\registers[23][25] ), .B1(n1847), .B2(
        \registers[22][25] ), .ZN(n1592) );
  AOI22_X1 U1331 ( .A1(n1836), .A2(\registers[25][25] ), .B1(n1835), .B2(
        \registers[24][25] ), .ZN(n1593) );
  AOI22_X1 U1332 ( .A1(n1824), .A2(\registers[31][25] ), .B1(n1823), .B2(
        \registers[30][25] ), .ZN(n1594) );
  AOI22_X1 U1333 ( .A1(n1848), .A2(\registers[23][26] ), .B1(n1847), .B2(
        \registers[22][26] ), .ZN(n1609) );
  AOI22_X1 U1334 ( .A1(n1836), .A2(\registers[25][26] ), .B1(n1835), .B2(
        \registers[24][26] ), .ZN(n1610) );
  AOI22_X1 U1335 ( .A1(n1824), .A2(\registers[31][26] ), .B1(n1823), .B2(
        \registers[30][26] ), .ZN(n1611) );
  AOI22_X1 U1336 ( .A1(n1848), .A2(\registers[23][27] ), .B1(n1847), .B2(
        \registers[22][27] ), .ZN(n1626) );
  AOI22_X1 U1337 ( .A1(n1836), .A2(\registers[25][27] ), .B1(n1835), .B2(
        \registers[24][27] ), .ZN(n1627) );
  AOI22_X1 U1338 ( .A1(n1824), .A2(\registers[31][27] ), .B1(n1823), .B2(
        \registers[30][27] ), .ZN(n1628) );
  AOI22_X1 U1339 ( .A1(n1848), .A2(\registers[23][28] ), .B1(n1847), .B2(
        \registers[22][28] ), .ZN(n1643) );
  AOI22_X1 U1340 ( .A1(n1836), .A2(\registers[25][28] ), .B1(n1835), .B2(
        \registers[24][28] ), .ZN(n1644) );
  AOI22_X1 U1341 ( .A1(n1824), .A2(\registers[31][28] ), .B1(n1823), .B2(
        \registers[30][28] ), .ZN(n1645) );
  AOI22_X1 U1342 ( .A1(n1848), .A2(\registers[23][29] ), .B1(n1847), .B2(
        \registers[22][29] ), .ZN(n1660) );
  AOI22_X1 U1343 ( .A1(n1836), .A2(\registers[25][29] ), .B1(n1835), .B2(
        \registers[24][29] ), .ZN(n1661) );
  AOI22_X1 U1344 ( .A1(n1824), .A2(\registers[31][29] ), .B1(n1823), .B2(
        \registers[30][29] ), .ZN(n1662) );
  AOI22_X1 U1345 ( .A1(n1848), .A2(\registers[23][30] ), .B1(n1847), .B2(
        \registers[22][30] ), .ZN(n1677) );
  AOI22_X1 U1346 ( .A1(n1836), .A2(\registers[25][30] ), .B1(n1835), .B2(
        \registers[24][30] ), .ZN(n1678) );
  AOI22_X1 U1347 ( .A1(n1824), .A2(\registers[31][30] ), .B1(n1823), .B2(
        \registers[30][30] ), .ZN(n1679) );
  AOI22_X1 U1348 ( .A1(n1848), .A2(\registers[23][31] ), .B1(n1847), .B2(
        \registers[22][31] ), .ZN(n1698) );
  AOI22_X1 U1349 ( .A1(n1836), .A2(\registers[25][31] ), .B1(n1835), .B2(
        \registers[24][31] ), .ZN(n1701) );
  AOI22_X1 U1350 ( .A1(n1824), .A2(\registers[31][31] ), .B1(n1823), .B2(
        \registers[30][31] ), .ZN(n1704) );
  AOI22_X1 U1351 ( .A1(\registers[23][8] ), .A2(n1942), .B1(\registers[22][8] ), .B2(n1939), .ZN(n716) );
  AOI22_X1 U1352 ( .A1(\registers[25][8] ), .A2(n1930), .B1(\registers[24][8] ), .B2(n1927), .ZN(n717) );
  AOI22_X1 U1353 ( .A1(\registers[31][8] ), .A2(n1918), .B1(\registers[30][8] ), .B2(n1915), .ZN(n718) );
  AOI22_X1 U1354 ( .A1(\registers[23][9] ), .A2(n1942), .B1(\registers[22][9] ), .B2(n1939), .ZN(n733) );
  AOI22_X1 U1355 ( .A1(\registers[25][9] ), .A2(n1930), .B1(\registers[24][9] ), .B2(n1927), .ZN(n734) );
  AOI22_X1 U1356 ( .A1(\registers[31][9] ), .A2(n1918), .B1(\registers[30][9] ), .B2(n1915), .ZN(n735) );
  AOI22_X1 U1357 ( .A1(\registers[23][10] ), .A2(n1942), .B1(
        \registers[22][10] ), .B2(n1939), .ZN(n750) );
  AOI22_X1 U1358 ( .A1(\registers[25][10] ), .A2(n1930), .B1(
        \registers[24][10] ), .B2(n1927), .ZN(n751) );
  AOI22_X1 U1359 ( .A1(\registers[31][10] ), .A2(n1918), .B1(
        \registers[30][10] ), .B2(n1915), .ZN(n752) );
  AOI22_X1 U1360 ( .A1(\registers[23][11] ), .A2(n1942), .B1(
        \registers[22][11] ), .B2(n1939), .ZN(n767) );
  AOI22_X1 U1361 ( .A1(\registers[25][11] ), .A2(n1930), .B1(
        \registers[24][11] ), .B2(n1927), .ZN(n768) );
  AOI22_X1 U1362 ( .A1(\registers[31][11] ), .A2(n1918), .B1(
        \registers[30][11] ), .B2(n1915), .ZN(n769) );
  AOI22_X1 U1363 ( .A1(\registers[23][12] ), .A2(n1942), .B1(
        \registers[22][12] ), .B2(n1939), .ZN(n784) );
  AOI22_X1 U1364 ( .A1(\registers[25][12] ), .A2(n1930), .B1(
        \registers[24][12] ), .B2(n1927), .ZN(n785) );
  AOI22_X1 U1365 ( .A1(\registers[31][12] ), .A2(n1918), .B1(
        \registers[30][12] ), .B2(n1915), .ZN(n786) );
  AOI22_X1 U1366 ( .A1(\registers[23][13] ), .A2(n1942), .B1(
        \registers[22][13] ), .B2(n1939), .ZN(n801) );
  AOI22_X1 U1367 ( .A1(\registers[25][13] ), .A2(n1930), .B1(
        \registers[24][13] ), .B2(n1927), .ZN(n802) );
  AOI22_X1 U1368 ( .A1(\registers[31][13] ), .A2(n1918), .B1(
        \registers[30][13] ), .B2(n1915), .ZN(n803) );
  AOI22_X1 U1369 ( .A1(\registers[23][14] ), .A2(n1942), .B1(
        \registers[22][14] ), .B2(n1939), .ZN(n818) );
  AOI22_X1 U1370 ( .A1(\registers[25][14] ), .A2(n1930), .B1(
        \registers[24][14] ), .B2(n1927), .ZN(n819) );
  AOI22_X1 U1371 ( .A1(\registers[31][14] ), .A2(n1918), .B1(
        \registers[30][14] ), .B2(n1915), .ZN(n820) );
  AOI22_X1 U1372 ( .A1(\registers[23][15] ), .A2(n1942), .B1(
        \registers[22][15] ), .B2(n1939), .ZN(n835) );
  AOI22_X1 U1373 ( .A1(\registers[25][15] ), .A2(n1930), .B1(
        \registers[24][15] ), .B2(n1927), .ZN(n836) );
  AOI22_X1 U1374 ( .A1(\registers[31][15] ), .A2(n1918), .B1(
        \registers[30][15] ), .B2(n1915), .ZN(n837) );
  AOI22_X1 U1375 ( .A1(\registers[23][16] ), .A2(n1942), .B1(
        \registers[22][16] ), .B2(n1939), .ZN(n852) );
  AOI22_X1 U1376 ( .A1(\registers[25][16] ), .A2(n1930), .B1(
        \registers[24][16] ), .B2(n1927), .ZN(n853) );
  AOI22_X1 U1377 ( .A1(\registers[31][16] ), .A2(n1918), .B1(
        \registers[30][16] ), .B2(n1915), .ZN(n854) );
  AOI22_X1 U1378 ( .A1(\registers[23][17] ), .A2(n1942), .B1(
        \registers[22][17] ), .B2(n1939), .ZN(n869) );
  AOI22_X1 U1379 ( .A1(\registers[25][17] ), .A2(n1930), .B1(
        \registers[24][17] ), .B2(n1927), .ZN(n870) );
  AOI22_X1 U1380 ( .A1(\registers[31][17] ), .A2(n1918), .B1(
        \registers[30][17] ), .B2(n1915), .ZN(n871) );
  AOI22_X1 U1381 ( .A1(\registers[23][18] ), .A2(n1942), .B1(
        \registers[22][18] ), .B2(n1939), .ZN(n886) );
  AOI22_X1 U1382 ( .A1(\registers[25][18] ), .A2(n1930), .B1(
        \registers[24][18] ), .B2(n1927), .ZN(n887) );
  AOI22_X1 U1383 ( .A1(\registers[31][18] ), .A2(n1918), .B1(
        \registers[30][18] ), .B2(n1915), .ZN(n888) );
  AOI22_X1 U1384 ( .A1(\registers[23][19] ), .A2(n1942), .B1(
        \registers[22][19] ), .B2(n1939), .ZN(n903) );
  AOI22_X1 U1385 ( .A1(\registers[25][19] ), .A2(n1930), .B1(
        \registers[24][19] ), .B2(n1927), .ZN(n904) );
  AOI22_X1 U1386 ( .A1(\registers[31][19] ), .A2(n1918), .B1(
        \registers[30][19] ), .B2(n1915), .ZN(n905) );
  AOI22_X1 U1387 ( .A1(\registers[23][20] ), .A2(n1941), .B1(
        \registers[22][20] ), .B2(n1938), .ZN(n920) );
  AOI22_X1 U1388 ( .A1(\registers[25][20] ), .A2(n1929), .B1(
        \registers[24][20] ), .B2(n1926), .ZN(n921) );
  AOI22_X1 U1389 ( .A1(\registers[31][20] ), .A2(n1917), .B1(
        \registers[30][20] ), .B2(n1914), .ZN(n922) );
  AOI22_X1 U1390 ( .A1(\registers[23][21] ), .A2(n1941), .B1(
        \registers[22][21] ), .B2(n1938), .ZN(n937) );
  AOI22_X1 U1391 ( .A1(\registers[25][21] ), .A2(n1929), .B1(
        \registers[24][21] ), .B2(n1926), .ZN(n938) );
  AOI22_X1 U1392 ( .A1(\registers[31][21] ), .A2(n1917), .B1(
        \registers[30][21] ), .B2(n1914), .ZN(n939) );
  AOI22_X1 U1393 ( .A1(\registers[23][22] ), .A2(n1941), .B1(
        \registers[22][22] ), .B2(n1938), .ZN(n954) );
  AOI22_X1 U1394 ( .A1(\registers[25][22] ), .A2(n1929), .B1(
        \registers[24][22] ), .B2(n1926), .ZN(n955) );
  AOI22_X1 U1395 ( .A1(\registers[31][22] ), .A2(n1917), .B1(
        \registers[30][22] ), .B2(n1914), .ZN(n956) );
  AOI22_X1 U1396 ( .A1(\registers[23][23] ), .A2(n1941), .B1(
        \registers[22][23] ), .B2(n1938), .ZN(n971) );
  AOI22_X1 U1397 ( .A1(\registers[25][23] ), .A2(n1929), .B1(
        \registers[24][23] ), .B2(n1926), .ZN(n972) );
  AOI22_X1 U1398 ( .A1(\registers[31][23] ), .A2(n1917), .B1(
        \registers[30][23] ), .B2(n1914), .ZN(n973) );
  AOI22_X1 U1399 ( .A1(\registers[23][24] ), .A2(n1941), .B1(
        \registers[22][24] ), .B2(n1938), .ZN(n988) );
  AOI22_X1 U1400 ( .A1(\registers[25][24] ), .A2(n1929), .B1(
        \registers[24][24] ), .B2(n1926), .ZN(n989) );
  AOI22_X1 U1401 ( .A1(\registers[31][24] ), .A2(n1917), .B1(
        \registers[30][24] ), .B2(n1914), .ZN(n990) );
  AOI22_X1 U1402 ( .A1(\registers[23][25] ), .A2(n1941), .B1(
        \registers[22][25] ), .B2(n1938), .ZN(n1005) );
  AOI22_X1 U1403 ( .A1(\registers[25][25] ), .A2(n1929), .B1(
        \registers[24][25] ), .B2(n1926), .ZN(n1006) );
  AOI22_X1 U1404 ( .A1(\registers[31][25] ), .A2(n1917), .B1(
        \registers[30][25] ), .B2(n1914), .ZN(n1007) );
  AOI22_X1 U1405 ( .A1(\registers[23][26] ), .A2(n1941), .B1(
        \registers[22][26] ), .B2(n1938), .ZN(n1022) );
  AOI22_X1 U1406 ( .A1(\registers[25][26] ), .A2(n1929), .B1(
        \registers[24][26] ), .B2(n1926), .ZN(n1023) );
  AOI22_X1 U1407 ( .A1(\registers[31][26] ), .A2(n1917), .B1(
        \registers[30][26] ), .B2(n1914), .ZN(n1024) );
  AOI22_X1 U1408 ( .A1(\registers[23][27] ), .A2(n1941), .B1(
        \registers[22][27] ), .B2(n1938), .ZN(n1039) );
  AOI22_X1 U1409 ( .A1(\registers[25][27] ), .A2(n1929), .B1(
        \registers[24][27] ), .B2(n1926), .ZN(n1040) );
  AOI22_X1 U1410 ( .A1(\registers[31][27] ), .A2(n1917), .B1(
        \registers[30][27] ), .B2(n1914), .ZN(n1041) );
  AOI22_X1 U1411 ( .A1(\registers[23][28] ), .A2(n1941), .B1(
        \registers[22][28] ), .B2(n1938), .ZN(n1056) );
  AOI22_X1 U1412 ( .A1(\registers[25][28] ), .A2(n1929), .B1(
        \registers[24][28] ), .B2(n1926), .ZN(n1057) );
  AOI22_X1 U1413 ( .A1(\registers[31][28] ), .A2(n1917), .B1(
        \registers[30][28] ), .B2(n1914), .ZN(n1058) );
  AOI22_X1 U1414 ( .A1(\registers[23][29] ), .A2(n1941), .B1(
        \registers[22][29] ), .B2(n1938), .ZN(n1073) );
  AOI22_X1 U1415 ( .A1(\registers[25][29] ), .A2(n1929), .B1(
        \registers[24][29] ), .B2(n1926), .ZN(n1074) );
  AOI22_X1 U1416 ( .A1(\registers[31][29] ), .A2(n1917), .B1(
        \registers[30][29] ), .B2(n1914), .ZN(n1075) );
  AOI22_X1 U1417 ( .A1(\registers[23][30] ), .A2(n1941), .B1(
        \registers[22][30] ), .B2(n1938), .ZN(n1090) );
  AOI22_X1 U1418 ( .A1(\registers[25][30] ), .A2(n1929), .B1(
        \registers[24][30] ), .B2(n1926), .ZN(n1091) );
  AOI22_X1 U1419 ( .A1(\registers[31][30] ), .A2(n1917), .B1(
        \registers[30][30] ), .B2(n1914), .ZN(n1092) );
  AOI22_X1 U1420 ( .A1(\registers[23][31] ), .A2(n1941), .B1(
        \registers[22][31] ), .B2(n1938), .ZN(n1111) );
  AOI22_X1 U1421 ( .A1(\registers[25][31] ), .A2(n1929), .B1(
        \registers[24][31] ), .B2(n1926), .ZN(n1114) );
  AOI22_X1 U1422 ( .A1(\registers[31][31] ), .A2(n1917), .B1(
        \registers[30][31] ), .B2(n1914), .ZN(n1117) );
  AND3_X1 U1423 ( .A1(add_rd1[3]), .A2(add_rd1[0]), .A3(add_rd1[4]), .ZN(n1703) );
  AND3_X1 U1424 ( .A1(add_rd1[3]), .A2(n2684), .A3(add_rd1[4]), .ZN(n1702) );
  AND3_X1 U1425 ( .A1(add_rd2[3]), .A2(add_rd2[0]), .A3(add_rd2[4]), .ZN(n1116) );
  AND3_X1 U1426 ( .A1(n2684), .A2(n2681), .A3(add_rd1[4]), .ZN(n1694) );
  AND3_X1 U1427 ( .A1(add_rd1[0]), .A2(n2681), .A3(add_rd1[4]), .ZN(n1696) );
  AND3_X1 U1428 ( .A1(add_rd2[3]), .A2(n2688), .A3(add_rd2[4]), .ZN(n1115) );
  AND3_X1 U1429 ( .A1(add_rd2[0]), .A2(n2685), .A3(add_rd2[4]), .ZN(n1109) );
  AND3_X1 U1430 ( .A1(n2688), .A2(n2685), .A3(add_rd2[4]), .ZN(n1107) );
  INV_X1 U1431 ( .A(add_rd2[3]), .ZN(n2685) );
  INV_X1 U1432 ( .A(add_rd2[0]), .ZN(n2688) );
  NAND4_X1 U1433 ( .A1(n540), .A2(n541), .A3(n542), .A4(n543), .ZN(N274) );
  AOI211_X1 U1434 ( .C1(\registers[5][0] ), .C2(n1913), .A(n569), .B(n570), 
        .ZN(n542) );
  AOI221_X1 U1435 ( .B1(\registers[13][0] ), .B2(n1880), .C1(\registers[2][0] ), .C2(n1877), .A(n585), .ZN(n540) );
  AOI221_X1 U1436 ( .B1(\registers[15][0] ), .B2(n1892), .C1(
        \registers[12][0] ), .C2(n1889), .A(n580), .ZN(n541) );
  NAND4_X1 U1437 ( .A1(n588), .A2(n589), .A3(n590), .A4(n591), .ZN(N273) );
  AOI211_X1 U1438 ( .C1(\registers[5][1] ), .C2(n1913), .A(n600), .B(n601), 
        .ZN(n590) );
  AOI221_X1 U1439 ( .B1(\registers[13][1] ), .B2(n1880), .C1(\registers[2][1] ), .C2(n1877), .A(n604), .ZN(n588) );
  AOI221_X1 U1440 ( .B1(\registers[15][1] ), .B2(n1892), .C1(
        \registers[12][1] ), .C2(n1889), .A(n603), .ZN(n589) );
  NAND4_X1 U1441 ( .A1(n605), .A2(n606), .A3(n607), .A4(n608), .ZN(N272) );
  AOI211_X1 U1442 ( .C1(\registers[5][2] ), .C2(n1913), .A(n617), .B(n618), 
        .ZN(n607) );
  AOI221_X1 U1443 ( .B1(\registers[13][2] ), .B2(n1880), .C1(\registers[2][2] ), .C2(n1877), .A(n621), .ZN(n605) );
  AOI221_X1 U1444 ( .B1(\registers[15][2] ), .B2(n1892), .C1(
        \registers[12][2] ), .C2(n1889), .A(n620), .ZN(n606) );
  NAND4_X1 U1445 ( .A1(n622), .A2(n623), .A3(n624), .A4(n625), .ZN(N271) );
  AOI211_X1 U1446 ( .C1(\registers[5][3] ), .C2(n1913), .A(n634), .B(n635), 
        .ZN(n624) );
  AOI221_X1 U1447 ( .B1(\registers[13][3] ), .B2(n1880), .C1(\registers[2][3] ), .C2(n1877), .A(n638), .ZN(n622) );
  AOI221_X1 U1448 ( .B1(\registers[15][3] ), .B2(n1892), .C1(
        \registers[12][3] ), .C2(n1889), .A(n637), .ZN(n623) );
  NAND4_X1 U1449 ( .A1(n639), .A2(n640), .A3(n641), .A4(n642), .ZN(N270) );
  AOI211_X1 U1450 ( .C1(\registers[5][4] ), .C2(n1913), .A(n651), .B(n652), 
        .ZN(n641) );
  AOI221_X1 U1451 ( .B1(\registers[13][4] ), .B2(n1880), .C1(\registers[2][4] ), .C2(n1877), .A(n655), .ZN(n639) );
  AOI221_X1 U1452 ( .B1(\registers[15][4] ), .B2(n1892), .C1(
        \registers[12][4] ), .C2(n1889), .A(n654), .ZN(n640) );
  NAND4_X1 U1453 ( .A1(n656), .A2(n657), .A3(n658), .A4(n659), .ZN(N269) );
  AOI211_X1 U1454 ( .C1(\registers[5][5] ), .C2(n1913), .A(n668), .B(n669), 
        .ZN(n658) );
  AOI221_X1 U1455 ( .B1(\registers[13][5] ), .B2(n1880), .C1(\registers[2][5] ), .C2(n1877), .A(n672), .ZN(n656) );
  AOI221_X1 U1456 ( .B1(\registers[15][5] ), .B2(n1892), .C1(
        \registers[12][5] ), .C2(n1889), .A(n671), .ZN(n657) );
  NAND4_X1 U1457 ( .A1(n673), .A2(n674), .A3(n675), .A4(n676), .ZN(N268) );
  AOI211_X1 U1458 ( .C1(\registers[5][6] ), .C2(n1913), .A(n685), .B(n686), 
        .ZN(n675) );
  AOI221_X1 U1459 ( .B1(\registers[13][6] ), .B2(n1880), .C1(\registers[2][6] ), .C2(n1877), .A(n689), .ZN(n673) );
  AOI221_X1 U1460 ( .B1(\registers[15][6] ), .B2(n1892), .C1(
        \registers[12][6] ), .C2(n1889), .A(n688), .ZN(n674) );
  NAND4_X1 U1461 ( .A1(n690), .A2(n691), .A3(n692), .A4(n693), .ZN(N267) );
  AOI211_X1 U1462 ( .C1(\registers[5][7] ), .C2(n1913), .A(n702), .B(n703), 
        .ZN(n692) );
  AOI221_X1 U1463 ( .B1(\registers[13][7] ), .B2(n1880), .C1(\registers[2][7] ), .C2(n1877), .A(n706), .ZN(n690) );
  AOI221_X1 U1464 ( .B1(\registers[15][7] ), .B2(n1892), .C1(
        \registers[12][7] ), .C2(n1889), .A(n705), .ZN(n691) );
  NAND4_X1 U1465 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(N177)
         );
  AOI211_X1 U1466 ( .C1(n1820), .C2(\registers[5][0] ), .A(n1156), .B(n1157), 
        .ZN(n1129) );
  AOI221_X1 U1467 ( .B1(n1787), .B2(\registers[13][0] ), .C1(n1784), .C2(
        \registers[2][0] ), .A(n1172), .ZN(n1127) );
  AOI221_X1 U1468 ( .B1(n1799), .B2(\registers[15][0] ), .C1(n1796), .C2(
        \registers[12][0] ), .A(n1167), .ZN(n1128) );
  NAND4_X1 U1469 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(N176)
         );
  AOI211_X1 U1470 ( .C1(n1820), .C2(\registers[5][1] ), .A(n1187), .B(n1188), 
        .ZN(n1177) );
  AOI221_X1 U1471 ( .B1(n1787), .B2(\registers[13][1] ), .C1(n1784), .C2(
        \registers[2][1] ), .A(n1191), .ZN(n1175) );
  AOI221_X1 U1472 ( .B1(n1799), .B2(\registers[15][1] ), .C1(n1796), .C2(
        \registers[12][1] ), .A(n1190), .ZN(n1176) );
  NAND4_X1 U1473 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(N175)
         );
  AOI211_X1 U1474 ( .C1(n1820), .C2(\registers[5][2] ), .A(n1204), .B(n1205), 
        .ZN(n1194) );
  AOI221_X1 U1475 ( .B1(n1787), .B2(\registers[13][2] ), .C1(n1784), .C2(
        \registers[2][2] ), .A(n1208), .ZN(n1192) );
  AOI221_X1 U1476 ( .B1(n1799), .B2(\registers[15][2] ), .C1(n1796), .C2(
        \registers[12][2] ), .A(n1207), .ZN(n1193) );
  NAND4_X1 U1477 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(N174)
         );
  AOI211_X1 U1478 ( .C1(n1820), .C2(\registers[5][3] ), .A(n1221), .B(n1222), 
        .ZN(n1211) );
  AOI221_X1 U1479 ( .B1(n1787), .B2(\registers[13][3] ), .C1(n1784), .C2(
        \registers[2][3] ), .A(n1225), .ZN(n1209) );
  AOI221_X1 U1480 ( .B1(n1799), .B2(\registers[15][3] ), .C1(n1796), .C2(
        \registers[12][3] ), .A(n1224), .ZN(n1210) );
  NAND4_X1 U1481 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(N173)
         );
  AOI211_X1 U1482 ( .C1(n1820), .C2(\registers[5][4] ), .A(n1238), .B(n1239), 
        .ZN(n1228) );
  AOI221_X1 U1483 ( .B1(n1787), .B2(\registers[13][4] ), .C1(n1784), .C2(
        \registers[2][4] ), .A(n1242), .ZN(n1226) );
  AOI221_X1 U1484 ( .B1(n1799), .B2(\registers[15][4] ), .C1(n1796), .C2(
        \registers[12][4] ), .A(n1241), .ZN(n1227) );
  NAND4_X1 U1485 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(N172)
         );
  AOI211_X1 U1486 ( .C1(n1820), .C2(\registers[5][5] ), .A(n1255), .B(n1256), 
        .ZN(n1245) );
  AOI221_X1 U1487 ( .B1(n1787), .B2(\registers[13][5] ), .C1(n1784), .C2(
        \registers[2][5] ), .A(n1259), .ZN(n1243) );
  AOI221_X1 U1488 ( .B1(n1799), .B2(\registers[15][5] ), .C1(n1796), .C2(
        \registers[12][5] ), .A(n1258), .ZN(n1244) );
  NAND4_X1 U1489 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(N171)
         );
  AOI211_X1 U1490 ( .C1(n1820), .C2(\registers[5][6] ), .A(n1272), .B(n1273), 
        .ZN(n1262) );
  AOI221_X1 U1491 ( .B1(n1787), .B2(\registers[13][6] ), .C1(n1784), .C2(
        \registers[2][6] ), .A(n1276), .ZN(n1260) );
  AOI221_X1 U1492 ( .B1(n1799), .B2(\registers[15][6] ), .C1(n1796), .C2(
        \registers[12][6] ), .A(n1275), .ZN(n1261) );
  NAND4_X1 U1493 ( .A1(n1277), .A2(n1278), .A3(n1279), .A4(n1280), .ZN(N170)
         );
  AOI211_X1 U1494 ( .C1(n1820), .C2(\registers[5][7] ), .A(n1289), .B(n1290), 
        .ZN(n1279) );
  AOI221_X1 U1495 ( .B1(n1787), .B2(\registers[13][7] ), .C1(n1784), .C2(
        \registers[2][7] ), .A(n1293), .ZN(n1277) );
  AOI221_X1 U1496 ( .B1(n1799), .B2(\registers[15][7] ), .C1(n1796), .C2(
        \registers[12][7] ), .A(n1292), .ZN(n1278) );
  NAND4_X1 U1497 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(N169)
         );
  AOI211_X1 U1498 ( .C1(n1819), .C2(\registers[5][8] ), .A(n1306), .B(n1307), 
        .ZN(n1296) );
  AOI221_X1 U1499 ( .B1(n1786), .B2(\registers[13][8] ), .C1(n1783), .C2(
        \registers[2][8] ), .A(n1310), .ZN(n1294) );
  AOI221_X1 U1500 ( .B1(n1798), .B2(\registers[15][8] ), .C1(n1795), .C2(
        \registers[12][8] ), .A(n1309), .ZN(n1295) );
  NAND4_X1 U1501 ( .A1(n1311), .A2(n1312), .A3(n1313), .A4(n1314), .ZN(N168)
         );
  AOI211_X1 U1502 ( .C1(n1819), .C2(\registers[5][9] ), .A(n1323), .B(n1324), 
        .ZN(n1313) );
  AOI221_X1 U1503 ( .B1(n1786), .B2(\registers[13][9] ), .C1(n1783), .C2(
        \registers[2][9] ), .A(n1327), .ZN(n1311) );
  AOI221_X1 U1504 ( .B1(n1798), .B2(\registers[15][9] ), .C1(n1795), .C2(
        \registers[12][9] ), .A(n1326), .ZN(n1312) );
  NAND4_X1 U1505 ( .A1(n1328), .A2(n1329), .A3(n1330), .A4(n1331), .ZN(N167)
         );
  AOI211_X1 U1506 ( .C1(n1819), .C2(\registers[5][10] ), .A(n1340), .B(n1341), 
        .ZN(n1330) );
  AOI221_X1 U1507 ( .B1(n1786), .B2(\registers[13][10] ), .C1(n1783), .C2(
        \registers[2][10] ), .A(n1344), .ZN(n1328) );
  AOI221_X1 U1508 ( .B1(n1798), .B2(\registers[15][10] ), .C1(n1795), .C2(
        \registers[12][10] ), .A(n1343), .ZN(n1329) );
  NAND4_X1 U1509 ( .A1(n1345), .A2(n1346), .A3(n1347), .A4(n1348), .ZN(N166)
         );
  AOI211_X1 U1510 ( .C1(n1819), .C2(\registers[5][11] ), .A(n1357), .B(n1358), 
        .ZN(n1347) );
  AOI221_X1 U1511 ( .B1(n1786), .B2(\registers[13][11] ), .C1(n1783), .C2(
        \registers[2][11] ), .A(n1361), .ZN(n1345) );
  AOI221_X1 U1512 ( .B1(n1798), .B2(\registers[15][11] ), .C1(n1795), .C2(
        \registers[12][11] ), .A(n1360), .ZN(n1346) );
  NAND4_X1 U1513 ( .A1(n1362), .A2(n1363), .A3(n1364), .A4(n1365), .ZN(N165)
         );
  AOI211_X1 U1514 ( .C1(n1819), .C2(\registers[5][12] ), .A(n1374), .B(n1375), 
        .ZN(n1364) );
  AOI221_X1 U1515 ( .B1(n1786), .B2(\registers[13][12] ), .C1(n1783), .C2(
        \registers[2][12] ), .A(n1378), .ZN(n1362) );
  AOI221_X1 U1516 ( .B1(n1798), .B2(\registers[15][12] ), .C1(n1795), .C2(
        \registers[12][12] ), .A(n1377), .ZN(n1363) );
  NAND4_X1 U1517 ( .A1(n1379), .A2(n1380), .A3(n1381), .A4(n1382), .ZN(N164)
         );
  AOI211_X1 U1518 ( .C1(n1819), .C2(\registers[5][13] ), .A(n1391), .B(n1392), 
        .ZN(n1381) );
  AOI221_X1 U1519 ( .B1(n1786), .B2(\registers[13][13] ), .C1(n1783), .C2(
        \registers[2][13] ), .A(n1395), .ZN(n1379) );
  AOI221_X1 U1520 ( .B1(n1798), .B2(\registers[15][13] ), .C1(n1795), .C2(
        \registers[12][13] ), .A(n1394), .ZN(n1380) );
  NAND4_X1 U1521 ( .A1(n1396), .A2(n1397), .A3(n1398), .A4(n1399), .ZN(N163)
         );
  AOI211_X1 U1522 ( .C1(n1819), .C2(\registers[5][14] ), .A(n1408), .B(n1409), 
        .ZN(n1398) );
  AOI221_X1 U1523 ( .B1(n1786), .B2(\registers[13][14] ), .C1(n1783), .C2(
        \registers[2][14] ), .A(n1412), .ZN(n1396) );
  AOI221_X1 U1524 ( .B1(n1798), .B2(\registers[15][14] ), .C1(n1795), .C2(
        \registers[12][14] ), .A(n1411), .ZN(n1397) );
  NAND4_X1 U1525 ( .A1(n1413), .A2(n1414), .A3(n1415), .A4(n1416), .ZN(N162)
         );
  AOI211_X1 U1526 ( .C1(n1819), .C2(\registers[5][15] ), .A(n1425), .B(n1426), 
        .ZN(n1415) );
  AOI221_X1 U1527 ( .B1(n1786), .B2(\registers[13][15] ), .C1(n1783), .C2(
        \registers[2][15] ), .A(n1429), .ZN(n1413) );
  AOI221_X1 U1528 ( .B1(n1798), .B2(\registers[15][15] ), .C1(n1795), .C2(
        \registers[12][15] ), .A(n1428), .ZN(n1414) );
  NAND4_X1 U1529 ( .A1(n1430), .A2(n1431), .A3(n1432), .A4(n1433), .ZN(N161)
         );
  AOI211_X1 U1530 ( .C1(n1819), .C2(\registers[5][16] ), .A(n1442), .B(n1443), 
        .ZN(n1432) );
  AOI221_X1 U1531 ( .B1(n1786), .B2(\registers[13][16] ), .C1(n1783), .C2(
        \registers[2][16] ), .A(n1446), .ZN(n1430) );
  AOI221_X1 U1532 ( .B1(n1798), .B2(\registers[15][16] ), .C1(n1795), .C2(
        \registers[12][16] ), .A(n1445), .ZN(n1431) );
  NAND4_X1 U1533 ( .A1(n1447), .A2(n1448), .A3(n1449), .A4(n1450), .ZN(N160)
         );
  AOI211_X1 U1534 ( .C1(n1819), .C2(\registers[5][17] ), .A(n1459), .B(n1460), 
        .ZN(n1449) );
  AOI221_X1 U1535 ( .B1(n1786), .B2(\registers[13][17] ), .C1(n1783), .C2(
        \registers[2][17] ), .A(n1463), .ZN(n1447) );
  AOI221_X1 U1536 ( .B1(n1798), .B2(\registers[15][17] ), .C1(n1795), .C2(
        \registers[12][17] ), .A(n1462), .ZN(n1448) );
  NAND4_X1 U1537 ( .A1(n1464), .A2(n1465), .A3(n1466), .A4(n1467), .ZN(N159)
         );
  AOI211_X1 U1538 ( .C1(n1819), .C2(\registers[5][18] ), .A(n1476), .B(n1477), 
        .ZN(n1466) );
  AOI221_X1 U1539 ( .B1(n1786), .B2(\registers[13][18] ), .C1(n1783), .C2(
        \registers[2][18] ), .A(n1480), .ZN(n1464) );
  AOI221_X1 U1540 ( .B1(n1798), .B2(\registers[15][18] ), .C1(n1795), .C2(
        \registers[12][18] ), .A(n1479), .ZN(n1465) );
  NAND4_X1 U1541 ( .A1(n1481), .A2(n1482), .A3(n1483), .A4(n1484), .ZN(N158)
         );
  AOI211_X1 U1542 ( .C1(n1819), .C2(\registers[5][19] ), .A(n1493), .B(n1494), 
        .ZN(n1483) );
  AOI221_X1 U1543 ( .B1(n1786), .B2(\registers[13][19] ), .C1(n1783), .C2(
        \registers[2][19] ), .A(n1497), .ZN(n1481) );
  AOI221_X1 U1544 ( .B1(n1798), .B2(\registers[15][19] ), .C1(n1795), .C2(
        \registers[12][19] ), .A(n1496), .ZN(n1482) );
  NAND4_X1 U1545 ( .A1(n1498), .A2(n1499), .A3(n1500), .A4(n1501), .ZN(N157)
         );
  AOI211_X1 U1546 ( .C1(n1818), .C2(\registers[5][20] ), .A(n1510), .B(n1511), 
        .ZN(n1500) );
  AOI221_X1 U1547 ( .B1(n1785), .B2(\registers[13][20] ), .C1(n1782), .C2(
        \registers[2][20] ), .A(n1514), .ZN(n1498) );
  AOI221_X1 U1548 ( .B1(n1797), .B2(\registers[15][20] ), .C1(n1794), .C2(
        \registers[12][20] ), .A(n1513), .ZN(n1499) );
  NAND4_X1 U1549 ( .A1(n1515), .A2(n1516), .A3(n1517), .A4(n1518), .ZN(N156)
         );
  AOI211_X1 U1550 ( .C1(n1818), .C2(\registers[5][21] ), .A(n1527), .B(n1528), 
        .ZN(n1517) );
  AOI221_X1 U1551 ( .B1(n1785), .B2(\registers[13][21] ), .C1(n1782), .C2(
        \registers[2][21] ), .A(n1531), .ZN(n1515) );
  AOI221_X1 U1552 ( .B1(n1797), .B2(\registers[15][21] ), .C1(n1794), .C2(
        \registers[12][21] ), .A(n1530), .ZN(n1516) );
  NAND4_X1 U1553 ( .A1(n1532), .A2(n1533), .A3(n1534), .A4(n1535), .ZN(N155)
         );
  AOI211_X1 U1554 ( .C1(n1818), .C2(\registers[5][22] ), .A(n1544), .B(n1545), 
        .ZN(n1534) );
  AOI221_X1 U1555 ( .B1(n1785), .B2(\registers[13][22] ), .C1(n1782), .C2(
        \registers[2][22] ), .A(n1548), .ZN(n1532) );
  AOI221_X1 U1556 ( .B1(n1797), .B2(\registers[15][22] ), .C1(n1794), .C2(
        \registers[12][22] ), .A(n1547), .ZN(n1533) );
  NAND4_X1 U1557 ( .A1(n1549), .A2(n1550), .A3(n1551), .A4(n1552), .ZN(N154)
         );
  AOI211_X1 U1558 ( .C1(n1818), .C2(\registers[5][23] ), .A(n1561), .B(n1562), 
        .ZN(n1551) );
  AOI221_X1 U1559 ( .B1(n1785), .B2(\registers[13][23] ), .C1(n1782), .C2(
        \registers[2][23] ), .A(n1565), .ZN(n1549) );
  AOI221_X1 U1560 ( .B1(n1797), .B2(\registers[15][23] ), .C1(n1794), .C2(
        \registers[12][23] ), .A(n1564), .ZN(n1550) );
  NAND4_X1 U1561 ( .A1(n1566), .A2(n1567), .A3(n1568), .A4(n1569), .ZN(N153)
         );
  AOI211_X1 U1562 ( .C1(n1818), .C2(\registers[5][24] ), .A(n1578), .B(n1579), 
        .ZN(n1568) );
  AOI221_X1 U1563 ( .B1(n1785), .B2(\registers[13][24] ), .C1(n1782), .C2(
        \registers[2][24] ), .A(n1582), .ZN(n1566) );
  AOI221_X1 U1564 ( .B1(n1797), .B2(\registers[15][24] ), .C1(n1794), .C2(
        \registers[12][24] ), .A(n1581), .ZN(n1567) );
  NAND4_X1 U1565 ( .A1(n1583), .A2(n1584), .A3(n1585), .A4(n1586), .ZN(N152)
         );
  AOI211_X1 U1566 ( .C1(n1818), .C2(\registers[5][25] ), .A(n1595), .B(n1596), 
        .ZN(n1585) );
  AOI221_X1 U1567 ( .B1(n1785), .B2(\registers[13][25] ), .C1(n1782), .C2(
        \registers[2][25] ), .A(n1599), .ZN(n1583) );
  AOI221_X1 U1568 ( .B1(n1797), .B2(\registers[15][25] ), .C1(n1794), .C2(
        \registers[12][25] ), .A(n1598), .ZN(n1584) );
  NAND4_X1 U1569 ( .A1(n1600), .A2(n1601), .A3(n1602), .A4(n1603), .ZN(N151)
         );
  AOI211_X1 U1570 ( .C1(n1818), .C2(\registers[5][26] ), .A(n1612), .B(n1613), 
        .ZN(n1602) );
  AOI221_X1 U1571 ( .B1(n1785), .B2(\registers[13][26] ), .C1(n1782), .C2(
        \registers[2][26] ), .A(n1616), .ZN(n1600) );
  AOI221_X1 U1572 ( .B1(n1797), .B2(\registers[15][26] ), .C1(n1794), .C2(
        \registers[12][26] ), .A(n1615), .ZN(n1601) );
  NAND4_X1 U1573 ( .A1(n1617), .A2(n1618), .A3(n1619), .A4(n1620), .ZN(N150)
         );
  AOI211_X1 U1574 ( .C1(n1818), .C2(\registers[5][27] ), .A(n1629), .B(n1630), 
        .ZN(n1619) );
  AOI221_X1 U1575 ( .B1(n1785), .B2(\registers[13][27] ), .C1(n1782), .C2(
        \registers[2][27] ), .A(n1633), .ZN(n1617) );
  AOI221_X1 U1576 ( .B1(n1797), .B2(\registers[15][27] ), .C1(n1794), .C2(
        \registers[12][27] ), .A(n1632), .ZN(n1618) );
  NAND4_X1 U1577 ( .A1(n1634), .A2(n1635), .A3(n1636), .A4(n1637), .ZN(N149)
         );
  AOI211_X1 U1578 ( .C1(n1818), .C2(\registers[5][28] ), .A(n1646), .B(n1647), 
        .ZN(n1636) );
  AOI221_X1 U1579 ( .B1(n1785), .B2(\registers[13][28] ), .C1(n1782), .C2(
        \registers[2][28] ), .A(n1650), .ZN(n1634) );
  AOI221_X1 U1580 ( .B1(n1797), .B2(\registers[15][28] ), .C1(n1794), .C2(
        \registers[12][28] ), .A(n1649), .ZN(n1635) );
  NAND4_X1 U1581 ( .A1(n1651), .A2(n1652), .A3(n1653), .A4(n1654), .ZN(N148)
         );
  AOI211_X1 U1582 ( .C1(n1818), .C2(\registers[5][29] ), .A(n1663), .B(n1664), 
        .ZN(n1653) );
  AOI221_X1 U1583 ( .B1(n1785), .B2(\registers[13][29] ), .C1(n1782), .C2(
        \registers[2][29] ), .A(n1667), .ZN(n1651) );
  AOI221_X1 U1584 ( .B1(n1797), .B2(\registers[15][29] ), .C1(n1794), .C2(
        \registers[12][29] ), .A(n1666), .ZN(n1652) );
  NAND4_X1 U1585 ( .A1(n1668), .A2(n1669), .A3(n1670), .A4(n1671), .ZN(N147)
         );
  AOI211_X1 U1586 ( .C1(n1818), .C2(\registers[5][30] ), .A(n1680), .B(n1681), 
        .ZN(n1670) );
  AOI221_X1 U1587 ( .B1(n1785), .B2(\registers[13][30] ), .C1(n1782), .C2(
        \registers[2][30] ), .A(n1684), .ZN(n1668) );
  AOI221_X1 U1588 ( .B1(n1797), .B2(\registers[15][30] ), .C1(n1794), .C2(
        \registers[12][30] ), .A(n1683), .ZN(n1669) );
  NAND4_X1 U1589 ( .A1(n1685), .A2(n1686), .A3(n1687), .A4(n1688), .ZN(N146)
         );
  AOI211_X1 U1590 ( .C1(n1818), .C2(\registers[5][31] ), .A(n1705), .B(n1706), 
        .ZN(n1687) );
  AOI221_X1 U1591 ( .B1(n1785), .B2(\registers[13][31] ), .C1(n1782), .C2(
        \registers[2][31] ), .A(n1713), .ZN(n1685) );
  AOI221_X1 U1592 ( .B1(n1797), .B2(\registers[15][31] ), .C1(n1794), .C2(
        \registers[12][31] ), .A(n1711), .ZN(n1686) );
  NAND4_X1 U1593 ( .A1(n707), .A2(n708), .A3(n709), .A4(n710), .ZN(N266) );
  AOI211_X1 U1594 ( .C1(\registers[5][8] ), .C2(n1912), .A(n719), .B(n720), 
        .ZN(n709) );
  AOI221_X1 U1595 ( .B1(\registers[13][8] ), .B2(n1879), .C1(\registers[2][8] ), .C2(n1876), .A(n723), .ZN(n707) );
  AOI221_X1 U1596 ( .B1(\registers[15][8] ), .B2(n1891), .C1(
        \registers[12][8] ), .C2(n1888), .A(n722), .ZN(n708) );
  NAND4_X1 U1597 ( .A1(n724), .A2(n725), .A3(n726), .A4(n727), .ZN(N265) );
  AOI211_X1 U1598 ( .C1(\registers[5][9] ), .C2(n1912), .A(n736), .B(n737), 
        .ZN(n726) );
  AOI221_X1 U1599 ( .B1(\registers[13][9] ), .B2(n1879), .C1(\registers[2][9] ), .C2(n1876), .A(n740), .ZN(n724) );
  AOI221_X1 U1600 ( .B1(\registers[15][9] ), .B2(n1891), .C1(
        \registers[12][9] ), .C2(n1888), .A(n739), .ZN(n725) );
  NAND4_X1 U1601 ( .A1(n741), .A2(n742), .A3(n743), .A4(n744), .ZN(N264) );
  AOI211_X1 U1602 ( .C1(\registers[5][10] ), .C2(n1912), .A(n753), .B(n754), 
        .ZN(n743) );
  AOI221_X1 U1603 ( .B1(\registers[13][10] ), .B2(n1879), .C1(
        \registers[2][10] ), .C2(n1876), .A(n757), .ZN(n741) );
  AOI221_X1 U1604 ( .B1(\registers[15][10] ), .B2(n1891), .C1(
        \registers[12][10] ), .C2(n1888), .A(n756), .ZN(n742) );
  NAND4_X1 U1605 ( .A1(n758), .A2(n759), .A3(n760), .A4(n761), .ZN(N263) );
  AOI211_X1 U1606 ( .C1(\registers[5][11] ), .C2(n1912), .A(n770), .B(n771), 
        .ZN(n760) );
  AOI221_X1 U1607 ( .B1(\registers[13][11] ), .B2(n1879), .C1(
        \registers[2][11] ), .C2(n1876), .A(n774), .ZN(n758) );
  AOI221_X1 U1608 ( .B1(\registers[15][11] ), .B2(n1891), .C1(
        \registers[12][11] ), .C2(n1888), .A(n773), .ZN(n759) );
  NAND4_X1 U1609 ( .A1(n775), .A2(n776), .A3(n777), .A4(n778), .ZN(N262) );
  AOI211_X1 U1610 ( .C1(\registers[5][12] ), .C2(n1912), .A(n787), .B(n788), 
        .ZN(n777) );
  AOI221_X1 U1611 ( .B1(\registers[13][12] ), .B2(n1879), .C1(
        \registers[2][12] ), .C2(n1876), .A(n791), .ZN(n775) );
  AOI221_X1 U1612 ( .B1(\registers[15][12] ), .B2(n1891), .C1(
        \registers[12][12] ), .C2(n1888), .A(n790), .ZN(n776) );
  NAND4_X1 U1613 ( .A1(n792), .A2(n793), .A3(n794), .A4(n795), .ZN(N261) );
  AOI211_X1 U1614 ( .C1(\registers[5][13] ), .C2(n1912), .A(n804), .B(n805), 
        .ZN(n794) );
  AOI221_X1 U1615 ( .B1(\registers[13][13] ), .B2(n1879), .C1(
        \registers[2][13] ), .C2(n1876), .A(n808), .ZN(n792) );
  AOI221_X1 U1616 ( .B1(\registers[15][13] ), .B2(n1891), .C1(
        \registers[12][13] ), .C2(n1888), .A(n807), .ZN(n793) );
  NAND4_X1 U1617 ( .A1(n809), .A2(n810), .A3(n811), .A4(n812), .ZN(N260) );
  AOI211_X1 U1618 ( .C1(\registers[5][14] ), .C2(n1912), .A(n821), .B(n822), 
        .ZN(n811) );
  AOI221_X1 U1619 ( .B1(\registers[13][14] ), .B2(n1879), .C1(
        \registers[2][14] ), .C2(n1876), .A(n825), .ZN(n809) );
  AOI221_X1 U1620 ( .B1(\registers[15][14] ), .B2(n1891), .C1(
        \registers[12][14] ), .C2(n1888), .A(n824), .ZN(n810) );
  NAND4_X1 U1621 ( .A1(n826), .A2(n827), .A3(n828), .A4(n829), .ZN(N259) );
  AOI211_X1 U1622 ( .C1(\registers[5][15] ), .C2(n1912), .A(n838), .B(n839), 
        .ZN(n828) );
  AOI221_X1 U1623 ( .B1(\registers[13][15] ), .B2(n1879), .C1(
        \registers[2][15] ), .C2(n1876), .A(n842), .ZN(n826) );
  AOI221_X1 U1624 ( .B1(\registers[15][15] ), .B2(n1891), .C1(
        \registers[12][15] ), .C2(n1888), .A(n841), .ZN(n827) );
  NAND4_X1 U1625 ( .A1(n843), .A2(n844), .A3(n845), .A4(n846), .ZN(N258) );
  AOI211_X1 U1626 ( .C1(\registers[5][16] ), .C2(n1912), .A(n855), .B(n856), 
        .ZN(n845) );
  AOI221_X1 U1627 ( .B1(\registers[13][16] ), .B2(n1879), .C1(
        \registers[2][16] ), .C2(n1876), .A(n859), .ZN(n843) );
  AOI221_X1 U1628 ( .B1(\registers[15][16] ), .B2(n1891), .C1(
        \registers[12][16] ), .C2(n1888), .A(n858), .ZN(n844) );
  NAND4_X1 U1629 ( .A1(n860), .A2(n861), .A3(n862), .A4(n863), .ZN(N257) );
  AOI211_X1 U1630 ( .C1(\registers[5][17] ), .C2(n1912), .A(n872), .B(n873), 
        .ZN(n862) );
  AOI221_X1 U1631 ( .B1(\registers[13][17] ), .B2(n1879), .C1(
        \registers[2][17] ), .C2(n1876), .A(n876), .ZN(n860) );
  AOI221_X1 U1632 ( .B1(\registers[15][17] ), .B2(n1891), .C1(
        \registers[12][17] ), .C2(n1888), .A(n875), .ZN(n861) );
  NAND4_X1 U1633 ( .A1(n877), .A2(n878), .A3(n879), .A4(n880), .ZN(N256) );
  AOI211_X1 U1634 ( .C1(\registers[5][18] ), .C2(n1912), .A(n889), .B(n890), 
        .ZN(n879) );
  AOI221_X1 U1635 ( .B1(\registers[13][18] ), .B2(n1879), .C1(
        \registers[2][18] ), .C2(n1876), .A(n893), .ZN(n877) );
  AOI221_X1 U1636 ( .B1(\registers[15][18] ), .B2(n1891), .C1(
        \registers[12][18] ), .C2(n1888), .A(n892), .ZN(n878) );
  NAND4_X1 U1637 ( .A1(n894), .A2(n895), .A3(n896), .A4(n897), .ZN(N255) );
  AOI211_X1 U1638 ( .C1(\registers[5][19] ), .C2(n1912), .A(n906), .B(n907), 
        .ZN(n896) );
  AOI221_X1 U1639 ( .B1(\registers[13][19] ), .B2(n1879), .C1(
        \registers[2][19] ), .C2(n1876), .A(n910), .ZN(n894) );
  AOI221_X1 U1640 ( .B1(\registers[15][19] ), .B2(n1891), .C1(
        \registers[12][19] ), .C2(n1888), .A(n909), .ZN(n895) );
  NAND4_X1 U1641 ( .A1(n911), .A2(n912), .A3(n913), .A4(n914), .ZN(N254) );
  AOI211_X1 U1642 ( .C1(\registers[5][20] ), .C2(n1911), .A(n923), .B(n924), 
        .ZN(n913) );
  AOI221_X1 U1643 ( .B1(\registers[13][20] ), .B2(n1878), .C1(
        \registers[2][20] ), .C2(n1875), .A(n927), .ZN(n911) );
  AOI221_X1 U1644 ( .B1(\registers[15][20] ), .B2(n1890), .C1(
        \registers[12][20] ), .C2(n1887), .A(n926), .ZN(n912) );
  NAND4_X1 U1645 ( .A1(n928), .A2(n929), .A3(n930), .A4(n931), .ZN(N253) );
  AOI211_X1 U1646 ( .C1(\registers[5][21] ), .C2(n1911), .A(n940), .B(n941), 
        .ZN(n930) );
  AOI221_X1 U1647 ( .B1(\registers[13][21] ), .B2(n1878), .C1(
        \registers[2][21] ), .C2(n1875), .A(n944), .ZN(n928) );
  AOI221_X1 U1648 ( .B1(\registers[15][21] ), .B2(n1890), .C1(
        \registers[12][21] ), .C2(n1887), .A(n943), .ZN(n929) );
  NAND4_X1 U1649 ( .A1(n945), .A2(n946), .A3(n947), .A4(n948), .ZN(N252) );
  AOI211_X1 U1650 ( .C1(\registers[5][22] ), .C2(n1911), .A(n957), .B(n958), 
        .ZN(n947) );
  AOI221_X1 U1651 ( .B1(\registers[13][22] ), .B2(n1878), .C1(
        \registers[2][22] ), .C2(n1875), .A(n961), .ZN(n945) );
  AOI221_X1 U1652 ( .B1(\registers[15][22] ), .B2(n1890), .C1(
        \registers[12][22] ), .C2(n1887), .A(n960), .ZN(n946) );
  NAND4_X1 U1653 ( .A1(n962), .A2(n963), .A3(n964), .A4(n965), .ZN(N251) );
  AOI211_X1 U1654 ( .C1(\registers[5][23] ), .C2(n1911), .A(n974), .B(n975), 
        .ZN(n964) );
  AOI221_X1 U1655 ( .B1(\registers[13][23] ), .B2(n1878), .C1(
        \registers[2][23] ), .C2(n1875), .A(n978), .ZN(n962) );
  AOI221_X1 U1656 ( .B1(\registers[15][23] ), .B2(n1890), .C1(
        \registers[12][23] ), .C2(n1887), .A(n977), .ZN(n963) );
  NAND4_X1 U1657 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(N250) );
  AOI211_X1 U1658 ( .C1(\registers[5][24] ), .C2(n1911), .A(n991), .B(n992), 
        .ZN(n981) );
  AOI221_X1 U1659 ( .B1(\registers[13][24] ), .B2(n1878), .C1(
        \registers[2][24] ), .C2(n1875), .A(n995), .ZN(n979) );
  AOI221_X1 U1660 ( .B1(\registers[15][24] ), .B2(n1890), .C1(
        \registers[12][24] ), .C2(n1887), .A(n994), .ZN(n980) );
  NAND4_X1 U1661 ( .A1(n996), .A2(n997), .A3(n998), .A4(n999), .ZN(N249) );
  AOI211_X1 U1662 ( .C1(\registers[5][25] ), .C2(n1911), .A(n1008), .B(n1009), 
        .ZN(n998) );
  AOI221_X1 U1663 ( .B1(\registers[13][25] ), .B2(n1878), .C1(
        \registers[2][25] ), .C2(n1875), .A(n1012), .ZN(n996) );
  AOI221_X1 U1664 ( .B1(\registers[15][25] ), .B2(n1890), .C1(
        \registers[12][25] ), .C2(n1887), .A(n1011), .ZN(n997) );
  NAND4_X1 U1665 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(N248)
         );
  AOI211_X1 U1666 ( .C1(\registers[5][26] ), .C2(n1911), .A(n1025), .B(n1026), 
        .ZN(n1015) );
  AOI221_X1 U1667 ( .B1(\registers[13][26] ), .B2(n1878), .C1(
        \registers[2][26] ), .C2(n1875), .A(n1029), .ZN(n1013) );
  AOI221_X1 U1668 ( .B1(\registers[15][26] ), .B2(n1890), .C1(
        \registers[12][26] ), .C2(n1887), .A(n1028), .ZN(n1014) );
  NAND4_X1 U1669 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(N247)
         );
  AOI211_X1 U1670 ( .C1(\registers[5][27] ), .C2(n1911), .A(n1042), .B(n1043), 
        .ZN(n1032) );
  AOI221_X1 U1671 ( .B1(\registers[13][27] ), .B2(n1878), .C1(
        \registers[2][27] ), .C2(n1875), .A(n1046), .ZN(n1030) );
  AOI221_X1 U1672 ( .B1(\registers[15][27] ), .B2(n1890), .C1(
        \registers[12][27] ), .C2(n1887), .A(n1045), .ZN(n1031) );
  NAND4_X1 U1673 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(N246)
         );
  AOI211_X1 U1674 ( .C1(\registers[5][28] ), .C2(n1911), .A(n1059), .B(n1060), 
        .ZN(n1049) );
  AOI221_X1 U1675 ( .B1(\registers[13][28] ), .B2(n1878), .C1(
        \registers[2][28] ), .C2(n1875), .A(n1063), .ZN(n1047) );
  AOI221_X1 U1676 ( .B1(\registers[15][28] ), .B2(n1890), .C1(
        \registers[12][28] ), .C2(n1887), .A(n1062), .ZN(n1048) );
  NAND4_X1 U1677 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(N245)
         );
  AOI211_X1 U1678 ( .C1(\registers[5][29] ), .C2(n1911), .A(n1076), .B(n1077), 
        .ZN(n1066) );
  AOI221_X1 U1679 ( .B1(\registers[13][29] ), .B2(n1878), .C1(
        \registers[2][29] ), .C2(n1875), .A(n1080), .ZN(n1064) );
  AOI221_X1 U1680 ( .B1(\registers[15][29] ), .B2(n1890), .C1(
        \registers[12][29] ), .C2(n1887), .A(n1079), .ZN(n1065) );
  NAND4_X1 U1681 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(N244)
         );
  AOI211_X1 U1682 ( .C1(\registers[5][30] ), .C2(n1911), .A(n1093), .B(n1094), 
        .ZN(n1083) );
  AOI221_X1 U1683 ( .B1(\registers[13][30] ), .B2(n1878), .C1(
        \registers[2][30] ), .C2(n1875), .A(n1097), .ZN(n1081) );
  AOI221_X1 U1684 ( .B1(\registers[15][30] ), .B2(n1890), .C1(
        \registers[12][30] ), .C2(n1887), .A(n1096), .ZN(n1082) );
  NAND4_X1 U1685 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(N243)
         );
  AOI211_X1 U1686 ( .C1(\registers[5][31] ), .C2(n1911), .A(n1118), .B(n1119), 
        .ZN(n1100) );
  AOI221_X1 U1687 ( .B1(\registers[13][31] ), .B2(n1878), .C1(
        \registers[2][31] ), .C2(n1875), .A(n1126), .ZN(n1098) );
  AOI221_X1 U1688 ( .B1(\registers[15][31] ), .B2(n1890), .C1(
        \registers[12][31] ), .C2(n1887), .A(n1124), .ZN(n1099) );
  INV_X1 U1689 ( .A(add_rd1[3]), .ZN(n2681) );
  INV_X1 U1690 ( .A(add_rd1[0]), .ZN(n2684) );
  INV_X1 U1691 ( .A(add_rd2[2]), .ZN(n2686) );
  INV_X1 U1692 ( .A(add_rd2[1]), .ZN(n2687) );
  INV_X1 U1693 ( .A(add_wr[2]), .ZN(n2166) );
  INV_X1 U1694 ( .A(add_wr[0]), .ZN(n2168) );
  INV_X1 U1695 ( .A(add_wr[1]), .ZN(n2167) );
  INV_X1 U1696 ( .A(add_rd1[2]), .ZN(n2682) );
  INV_X1 U1697 ( .A(add_rd1[1]), .ZN(n2683) );
  INV_X1 U1698 ( .A(\registers[19][0] ), .ZN(n2488) );
  INV_X1 U1699 ( .A(\registers[21][0] ), .ZN(n2552) );
  INV_X1 U1700 ( .A(\registers[27][0] ), .ZN(n2616) );
  INV_X1 U1701 ( .A(\registers[29][0] ), .ZN(n2680) );
  INV_X1 U1702 ( .A(\registers[1][0] ), .ZN(n2200) );
  INV_X1 U1703 ( .A(\registers[19][1] ), .ZN(n2487) );
  INV_X1 U1704 ( .A(\registers[21][1] ), .ZN(n2551) );
  INV_X1 U1705 ( .A(\registers[27][1] ), .ZN(n2615) );
  INV_X1 U1706 ( .A(\registers[29][1] ), .ZN(n2679) );
  INV_X1 U1707 ( .A(\registers[1][1] ), .ZN(n2199) );
  INV_X1 U1708 ( .A(\registers[19][2] ), .ZN(n2486) );
  INV_X1 U1709 ( .A(\registers[21][2] ), .ZN(n2550) );
  INV_X1 U1710 ( .A(\registers[27][2] ), .ZN(n2614) );
  INV_X1 U1711 ( .A(\registers[29][2] ), .ZN(n2678) );
  INV_X1 U1712 ( .A(\registers[1][2] ), .ZN(n2198) );
  INV_X1 U1713 ( .A(\registers[19][3] ), .ZN(n2485) );
  INV_X1 U1714 ( .A(\registers[21][3] ), .ZN(n2549) );
  INV_X1 U1715 ( .A(\registers[27][3] ), .ZN(n2613) );
  INV_X1 U1716 ( .A(\registers[29][3] ), .ZN(n2677) );
  INV_X1 U1717 ( .A(\registers[1][3] ), .ZN(n2197) );
  INV_X1 U1718 ( .A(\registers[19][4] ), .ZN(n2484) );
  INV_X1 U1719 ( .A(\registers[21][4] ), .ZN(n2548) );
  INV_X1 U1720 ( .A(\registers[27][4] ), .ZN(n2612) );
  INV_X1 U1721 ( .A(\registers[29][4] ), .ZN(n2676) );
  INV_X1 U1722 ( .A(\registers[1][4] ), .ZN(n2196) );
  INV_X1 U1723 ( .A(\registers[19][5] ), .ZN(n2483) );
  INV_X1 U1724 ( .A(\registers[21][5] ), .ZN(n2547) );
  INV_X1 U1725 ( .A(\registers[27][5] ), .ZN(n2611) );
  INV_X1 U1726 ( .A(\registers[29][5] ), .ZN(n2675) );
  INV_X1 U1727 ( .A(\registers[1][5] ), .ZN(n2195) );
  INV_X1 U1728 ( .A(\registers[19][6] ), .ZN(n2482) );
  INV_X1 U1729 ( .A(\registers[21][6] ), .ZN(n2546) );
  INV_X1 U1730 ( .A(\registers[27][6] ), .ZN(n2610) );
  INV_X1 U1731 ( .A(\registers[29][6] ), .ZN(n2674) );
  INV_X1 U1732 ( .A(\registers[1][6] ), .ZN(n2194) );
  INV_X1 U1733 ( .A(\registers[19][7] ), .ZN(n2481) );
  INV_X1 U1734 ( .A(\registers[21][7] ), .ZN(n2545) );
  INV_X1 U1735 ( .A(\registers[27][7] ), .ZN(n2609) );
  INV_X1 U1736 ( .A(\registers[29][7] ), .ZN(n2673) );
  INV_X1 U1737 ( .A(\registers[1][7] ), .ZN(n2193) );
  INV_X1 U1738 ( .A(\registers[19][8] ), .ZN(n2480) );
  INV_X1 U1739 ( .A(\registers[21][8] ), .ZN(n2544) );
  INV_X1 U1740 ( .A(\registers[27][8] ), .ZN(n2608) );
  INV_X1 U1741 ( .A(\registers[29][8] ), .ZN(n2672) );
  INV_X1 U1742 ( .A(\registers[1][8] ), .ZN(n2192) );
  INV_X1 U1743 ( .A(\registers[19][9] ), .ZN(n2479) );
  INV_X1 U1744 ( .A(\registers[21][9] ), .ZN(n2543) );
  INV_X1 U1745 ( .A(\registers[27][9] ), .ZN(n2607) );
  INV_X1 U1746 ( .A(\registers[29][9] ), .ZN(n2671) );
  INV_X1 U1747 ( .A(\registers[1][9] ), .ZN(n2191) );
  INV_X1 U1748 ( .A(\registers[19][10] ), .ZN(n2478) );
  INV_X1 U1749 ( .A(\registers[21][10] ), .ZN(n2542) );
  INV_X1 U1750 ( .A(\registers[27][10] ), .ZN(n2606) );
  INV_X1 U1751 ( .A(\registers[29][10] ), .ZN(n2670) );
  INV_X1 U1752 ( .A(\registers[1][10] ), .ZN(n2190) );
  INV_X1 U1753 ( .A(\registers[19][11] ), .ZN(n2477) );
  INV_X1 U1754 ( .A(\registers[21][11] ), .ZN(n2541) );
  INV_X1 U1755 ( .A(\registers[27][11] ), .ZN(n2605) );
  INV_X1 U1756 ( .A(\registers[29][11] ), .ZN(n2669) );
  INV_X1 U1757 ( .A(\registers[1][11] ), .ZN(n2189) );
  INV_X1 U1758 ( .A(\registers[19][12] ), .ZN(n2476) );
  INV_X1 U1759 ( .A(\registers[21][12] ), .ZN(n2540) );
  INV_X1 U1760 ( .A(\registers[27][12] ), .ZN(n2604) );
  INV_X1 U1761 ( .A(\registers[29][12] ), .ZN(n2668) );
  INV_X1 U1762 ( .A(\registers[1][12] ), .ZN(n2188) );
  INV_X1 U1763 ( .A(\registers[19][13] ), .ZN(n2475) );
  INV_X1 U1764 ( .A(\registers[21][13] ), .ZN(n2539) );
  INV_X1 U1765 ( .A(\registers[27][13] ), .ZN(n2603) );
  INV_X1 U1766 ( .A(\registers[29][13] ), .ZN(n2667) );
  INV_X1 U1767 ( .A(\registers[1][13] ), .ZN(n2187) );
  INV_X1 U1768 ( .A(\registers[19][14] ), .ZN(n2474) );
  INV_X1 U1769 ( .A(\registers[21][14] ), .ZN(n2538) );
  INV_X1 U1770 ( .A(\registers[27][14] ), .ZN(n2602) );
  INV_X1 U1771 ( .A(\registers[29][14] ), .ZN(n2666) );
  INV_X1 U1772 ( .A(\registers[1][14] ), .ZN(n2186) );
  INV_X1 U1773 ( .A(\registers[19][15] ), .ZN(n2473) );
  INV_X1 U1774 ( .A(\registers[21][15] ), .ZN(n2537) );
  INV_X1 U1775 ( .A(\registers[27][15] ), .ZN(n2601) );
  INV_X1 U1776 ( .A(\registers[29][15] ), .ZN(n2665) );
  INV_X1 U1777 ( .A(\registers[1][15] ), .ZN(n2185) );
  INV_X1 U1778 ( .A(\registers[19][16] ), .ZN(n2472) );
  INV_X1 U1779 ( .A(\registers[21][16] ), .ZN(n2536) );
  INV_X1 U1780 ( .A(\registers[27][16] ), .ZN(n2600) );
  INV_X1 U1781 ( .A(\registers[29][16] ), .ZN(n2664) );
  INV_X1 U1782 ( .A(\registers[1][16] ), .ZN(n2184) );
  INV_X1 U1783 ( .A(\registers[19][17] ), .ZN(n2471) );
  INV_X1 U1784 ( .A(\registers[21][17] ), .ZN(n2535) );
  INV_X1 U1785 ( .A(\registers[27][17] ), .ZN(n2599) );
  INV_X1 U1786 ( .A(\registers[29][17] ), .ZN(n2663) );
  INV_X1 U1787 ( .A(\registers[1][17] ), .ZN(n2183) );
  INV_X1 U1788 ( .A(\registers[19][18] ), .ZN(n2470) );
  INV_X1 U1789 ( .A(\registers[21][18] ), .ZN(n2534) );
  INV_X1 U1790 ( .A(\registers[27][18] ), .ZN(n2598) );
  INV_X1 U1791 ( .A(\registers[29][18] ), .ZN(n2662) );
  INV_X1 U1792 ( .A(\registers[1][18] ), .ZN(n2182) );
  INV_X1 U1793 ( .A(\registers[19][19] ), .ZN(n2469) );
  INV_X1 U1794 ( .A(\registers[21][19] ), .ZN(n2533) );
  INV_X1 U1795 ( .A(\registers[27][19] ), .ZN(n2597) );
  INV_X1 U1796 ( .A(\registers[29][19] ), .ZN(n2661) );
  INV_X1 U1797 ( .A(\registers[1][19] ), .ZN(n2181) );
  INV_X1 U1798 ( .A(\registers[19][20] ), .ZN(n2468) );
  INV_X1 U1799 ( .A(\registers[21][20] ), .ZN(n2532) );
  INV_X1 U1800 ( .A(\registers[27][20] ), .ZN(n2596) );
  INV_X1 U1801 ( .A(\registers[29][20] ), .ZN(n2660) );
  INV_X1 U1802 ( .A(\registers[1][20] ), .ZN(n2180) );
  INV_X1 U1803 ( .A(\registers[19][21] ), .ZN(n2467) );
  INV_X1 U1804 ( .A(\registers[21][21] ), .ZN(n2531) );
  INV_X1 U1805 ( .A(\registers[27][21] ), .ZN(n2595) );
  INV_X1 U1806 ( .A(\registers[29][21] ), .ZN(n2659) );
  INV_X1 U1807 ( .A(\registers[1][21] ), .ZN(n2179) );
  INV_X1 U1808 ( .A(\registers[19][22] ), .ZN(n2466) );
  INV_X1 U1809 ( .A(\registers[21][22] ), .ZN(n2530) );
  INV_X1 U1810 ( .A(\registers[27][22] ), .ZN(n2594) );
  INV_X1 U1811 ( .A(\registers[29][22] ), .ZN(n2658) );
  INV_X1 U1812 ( .A(\registers[1][22] ), .ZN(n2178) );
  INV_X1 U1813 ( .A(\registers[19][23] ), .ZN(n2465) );
  INV_X1 U1814 ( .A(\registers[21][23] ), .ZN(n2529) );
  INV_X1 U1815 ( .A(\registers[27][23] ), .ZN(n2593) );
  INV_X1 U1816 ( .A(\registers[29][23] ), .ZN(n2657) );
  INV_X1 U1817 ( .A(\registers[1][23] ), .ZN(n2177) );
  INV_X1 U1818 ( .A(\registers[19][24] ), .ZN(n2464) );
  INV_X1 U1819 ( .A(\registers[21][24] ), .ZN(n2528) );
  INV_X1 U1820 ( .A(\registers[27][24] ), .ZN(n2592) );
  INV_X1 U1821 ( .A(\registers[29][24] ), .ZN(n2656) );
  INV_X1 U1822 ( .A(\registers[1][24] ), .ZN(n2176) );
  INV_X1 U1823 ( .A(\registers[19][25] ), .ZN(n2463) );
  INV_X1 U1824 ( .A(\registers[21][25] ), .ZN(n2527) );
  INV_X1 U1825 ( .A(\registers[27][25] ), .ZN(n2591) );
  INV_X1 U1826 ( .A(\registers[29][25] ), .ZN(n2655) );
  INV_X1 U1827 ( .A(\registers[1][25] ), .ZN(n2175) );
  INV_X1 U1828 ( .A(\registers[19][26] ), .ZN(n2462) );
  INV_X1 U1829 ( .A(\registers[21][26] ), .ZN(n2526) );
  INV_X1 U1830 ( .A(\registers[27][26] ), .ZN(n2590) );
  INV_X1 U1831 ( .A(\registers[29][26] ), .ZN(n2654) );
  INV_X1 U1844 ( .A(\registers[1][26] ), .ZN(n2174) );
  INV_X1 U1845 ( .A(\registers[19][27] ), .ZN(n2461) );
  INV_X1 U1846 ( .A(\registers[21][27] ), .ZN(n2525) );
  INV_X1 U1847 ( .A(\registers[27][27] ), .ZN(n2589) );
  INV_X1 U1848 ( .A(\registers[29][27] ), .ZN(n2653) );
  INV_X1 U1849 ( .A(\registers[1][27] ), .ZN(n2173) );
  INV_X1 U1850 ( .A(\registers[19][28] ), .ZN(n2460) );
  INV_X1 U1851 ( .A(\registers[21][28] ), .ZN(n2524) );
  INV_X1 U1852 ( .A(\registers[27][28] ), .ZN(n2588) );
  INV_X1 U1853 ( .A(\registers[29][28] ), .ZN(n2652) );
  INV_X1 U1854 ( .A(\registers[1][28] ), .ZN(n2172) );
  INV_X1 U1855 ( .A(\registers[19][29] ), .ZN(n2459) );
  INV_X1 U1856 ( .A(\registers[21][29] ), .ZN(n2523) );
  INV_X1 U1857 ( .A(\registers[27][29] ), .ZN(n2587) );
  INV_X1 U1858 ( .A(\registers[29][29] ), .ZN(n2651) );
  INV_X1 U1859 ( .A(\registers[1][29] ), .ZN(n2171) );
  INV_X1 U1860 ( .A(\registers[19][30] ), .ZN(n2458) );
  INV_X1 U1861 ( .A(\registers[21][30] ), .ZN(n2522) );
  INV_X1 U1862 ( .A(\registers[27][30] ), .ZN(n2586) );
  INV_X1 U1863 ( .A(\registers[29][30] ), .ZN(n2650) );
  INV_X1 U1864 ( .A(\registers[1][30] ), .ZN(n2170) );
  INV_X1 U1865 ( .A(\registers[19][31] ), .ZN(n2457) );
  INV_X1 U1866 ( .A(\registers[21][31] ), .ZN(n2521) );
  INV_X1 U1867 ( .A(\registers[27][31] ), .ZN(n2585) );
  INV_X1 U1868 ( .A(\registers[29][31] ), .ZN(n2649) );
  INV_X1 U1869 ( .A(\registers[1][31] ), .ZN(n2169) );
  INV_X1 U1870 ( .A(\registers[11][0] ), .ZN(n2392) );
  INV_X1 U1871 ( .A(\registers[9][0] ), .ZN(n2328) );
  INV_X1 U1872 ( .A(\registers[10][0] ), .ZN(n2360) );
  INV_X1 U1873 ( .A(\registers[11][1] ), .ZN(n2391) );
  INV_X1 U1874 ( .A(\registers[9][1] ), .ZN(n2327) );
  INV_X1 U1875 ( .A(\registers[10][1] ), .ZN(n2359) );
  INV_X1 U1876 ( .A(\registers[11][2] ), .ZN(n2390) );
  INV_X1 U1877 ( .A(\registers[9][2] ), .ZN(n2326) );
  INV_X1 U1878 ( .A(\registers[10][2] ), .ZN(n2358) );
  INV_X1 U1879 ( .A(\registers[11][3] ), .ZN(n2389) );
  INV_X1 U1880 ( .A(\registers[9][3] ), .ZN(n2325) );
  INV_X1 U1881 ( .A(\registers[10][3] ), .ZN(n2357) );
  INV_X1 U1882 ( .A(\registers[11][4] ), .ZN(n2388) );
  INV_X1 U1883 ( .A(\registers[9][4] ), .ZN(n2324) );
  INV_X1 U1884 ( .A(\registers[10][4] ), .ZN(n2356) );
  INV_X1 U1885 ( .A(\registers[11][5] ), .ZN(n2387) );
  INV_X1 U1886 ( .A(\registers[9][5] ), .ZN(n2323) );
  INV_X1 U1887 ( .A(\registers[10][5] ), .ZN(n2355) );
  INV_X1 U1888 ( .A(\registers[11][6] ), .ZN(n2386) );
  INV_X1 U1889 ( .A(\registers[9][6] ), .ZN(n2322) );
  INV_X1 U1890 ( .A(\registers[10][6] ), .ZN(n2354) );
  INV_X1 U1891 ( .A(\registers[11][7] ), .ZN(n2385) );
  INV_X1 U1892 ( .A(\registers[9][7] ), .ZN(n2321) );
  INV_X1 U1893 ( .A(\registers[10][7] ), .ZN(n2353) );
  INV_X1 U1894 ( .A(\registers[11][8] ), .ZN(n2384) );
  INV_X1 U1895 ( .A(\registers[9][8] ), .ZN(n2320) );
  INV_X1 U1896 ( .A(\registers[10][8] ), .ZN(n2352) );
  INV_X1 U1897 ( .A(\registers[11][9] ), .ZN(n2383) );
  INV_X1 U1898 ( .A(\registers[9][9] ), .ZN(n2319) );
  INV_X1 U1899 ( .A(\registers[10][9] ), .ZN(n2351) );
  INV_X1 U1900 ( .A(\registers[11][10] ), .ZN(n2382) );
  INV_X1 U1901 ( .A(\registers[9][10] ), .ZN(n2318) );
  INV_X1 U1902 ( .A(\registers[10][10] ), .ZN(n2350) );
  INV_X1 U1903 ( .A(\registers[11][11] ), .ZN(n2381) );
  INV_X1 U1904 ( .A(\registers[9][11] ), .ZN(n2317) );
  INV_X1 U1905 ( .A(\registers[10][11] ), .ZN(n2349) );
  INV_X1 U1906 ( .A(\registers[11][12] ), .ZN(n2380) );
  INV_X1 U1907 ( .A(\registers[9][12] ), .ZN(n2316) );
  INV_X1 U1908 ( .A(\registers[10][12] ), .ZN(n2348) );
  INV_X1 U1909 ( .A(\registers[11][13] ), .ZN(n2379) );
  INV_X1 U1910 ( .A(\registers[9][13] ), .ZN(n2315) );
  INV_X1 U1911 ( .A(\registers[10][13] ), .ZN(n2347) );
  INV_X1 U1912 ( .A(\registers[11][14] ), .ZN(n2378) );
  INV_X1 U1913 ( .A(\registers[9][14] ), .ZN(n2314) );
  INV_X1 U1914 ( .A(\registers[10][14] ), .ZN(n2346) );
  INV_X1 U1915 ( .A(\registers[11][15] ), .ZN(n2377) );
  INV_X1 U1916 ( .A(\registers[9][15] ), .ZN(n2313) );
  INV_X1 U1917 ( .A(\registers[10][15] ), .ZN(n2345) );
  INV_X1 U1918 ( .A(\registers[11][16] ), .ZN(n2376) );
  INV_X1 U1919 ( .A(\registers[9][16] ), .ZN(n2312) );
  INV_X1 U1920 ( .A(\registers[10][16] ), .ZN(n2344) );
  INV_X1 U1921 ( .A(\registers[11][17] ), .ZN(n2375) );
  INV_X1 U1922 ( .A(\registers[9][17] ), .ZN(n2311) );
  INV_X1 U1923 ( .A(\registers[10][17] ), .ZN(n2343) );
  INV_X1 U1924 ( .A(\registers[11][18] ), .ZN(n2374) );
  INV_X1 U1925 ( .A(\registers[9][18] ), .ZN(n2310) );
  INV_X1 U1926 ( .A(\registers[10][18] ), .ZN(n2342) );
  INV_X1 U1927 ( .A(\registers[11][19] ), .ZN(n2373) );
  INV_X1 U1928 ( .A(\registers[9][19] ), .ZN(n2309) );
  INV_X1 U1929 ( .A(\registers[10][19] ), .ZN(n2341) );
  INV_X1 U1930 ( .A(\registers[11][20] ), .ZN(n2372) );
  INV_X1 U1931 ( .A(\registers[9][20] ), .ZN(n2308) );
  INV_X1 U1932 ( .A(\registers[10][20] ), .ZN(n2340) );
  INV_X1 U1933 ( .A(\registers[11][21] ), .ZN(n2371) );
  INV_X1 U1934 ( .A(\registers[9][21] ), .ZN(n2307) );
  INV_X1 U1935 ( .A(\registers[10][21] ), .ZN(n2339) );
  INV_X1 U1936 ( .A(\registers[11][22] ), .ZN(n2370) );
  INV_X1 U1937 ( .A(\registers[9][22] ), .ZN(n2306) );
  INV_X1 U1938 ( .A(\registers[10][22] ), .ZN(n2338) );
  INV_X1 U1939 ( .A(\registers[11][23] ), .ZN(n2369) );
  INV_X1 U1940 ( .A(\registers[9][23] ), .ZN(n2305) );
  INV_X1 U1941 ( .A(\registers[10][23] ), .ZN(n2337) );
  INV_X1 U1942 ( .A(\registers[11][24] ), .ZN(n2368) );
  INV_X1 U1943 ( .A(\registers[9][24] ), .ZN(n2304) );
  INV_X1 U1944 ( .A(\registers[10][24] ), .ZN(n2336) );
  INV_X1 U1945 ( .A(\registers[11][25] ), .ZN(n2367) );
  INV_X1 U1946 ( .A(\registers[9][25] ), .ZN(n2303) );
  INV_X1 U1947 ( .A(\registers[10][25] ), .ZN(n2335) );
  INV_X1 U1948 ( .A(\registers[11][26] ), .ZN(n2366) );
  INV_X1 U1949 ( .A(\registers[9][26] ), .ZN(n2302) );
  INV_X1 U1950 ( .A(\registers[10][26] ), .ZN(n2334) );
  INV_X1 U1951 ( .A(\registers[11][27] ), .ZN(n2365) );
  INV_X1 U1952 ( .A(\registers[9][27] ), .ZN(n2301) );
  INV_X1 U1953 ( .A(\registers[10][27] ), .ZN(n2333) );
  INV_X1 U1954 ( .A(\registers[11][28] ), .ZN(n2364) );
  INV_X1 U1955 ( .A(\registers[9][28] ), .ZN(n2300) );
  INV_X1 U1956 ( .A(\registers[10][28] ), .ZN(n2332) );
  INV_X1 U1957 ( .A(\registers[11][29] ), .ZN(n2363) );
  INV_X1 U1958 ( .A(\registers[9][29] ), .ZN(n2299) );
  INV_X1 U1959 ( .A(\registers[10][29] ), .ZN(n2331) );
  INV_X1 U1960 ( .A(\registers[11][30] ), .ZN(n2362) );
  INV_X1 U1961 ( .A(\registers[9][30] ), .ZN(n2298) );
  INV_X1 U1962 ( .A(\registers[10][30] ), .ZN(n2330) );
  INV_X1 U1963 ( .A(\registers[11][31] ), .ZN(n2361) );
  INV_X1 U1964 ( .A(\registers[9][31] ), .ZN(n2297) );
  INV_X1 U1965 ( .A(\registers[10][31] ), .ZN(n2329) );
  INV_X1 U1966 ( .A(\registers[8][0] ), .ZN(n2296) );
  INV_X1 U1967 ( .A(\registers[14][0] ), .ZN(n2424) );
  INV_X1 U1968 ( .A(\registers[4][0] ), .ZN(n2232) );
  INV_X1 U1969 ( .A(\registers[8][1] ), .ZN(n2295) );
  INV_X1 U1970 ( .A(\registers[14][1] ), .ZN(n2423) );
  INV_X1 U1971 ( .A(\registers[4][1] ), .ZN(n2231) );
  INV_X1 U1972 ( .A(\registers[8][2] ), .ZN(n2294) );
  INV_X1 U1973 ( .A(\registers[14][2] ), .ZN(n2422) );
  INV_X1 U1974 ( .A(\registers[4][2] ), .ZN(n2230) );
  INV_X1 U1975 ( .A(\registers[8][3] ), .ZN(n2293) );
  INV_X1 U1976 ( .A(\registers[14][3] ), .ZN(n2421) );
  INV_X1 U1977 ( .A(\registers[4][3] ), .ZN(n2229) );
  INV_X1 U1978 ( .A(\registers[8][4] ), .ZN(n2292) );
  INV_X1 U1979 ( .A(\registers[14][4] ), .ZN(n2420) );
  INV_X1 U1980 ( .A(\registers[4][4] ), .ZN(n2228) );
  INV_X1 U1981 ( .A(\registers[8][5] ), .ZN(n2291) );
  INV_X1 U1982 ( .A(\registers[14][5] ), .ZN(n2419) );
  INV_X1 U1983 ( .A(\registers[4][5] ), .ZN(n2227) );
  INV_X1 U1984 ( .A(\registers[8][6] ), .ZN(n2290) );
  INV_X1 U1985 ( .A(\registers[14][6] ), .ZN(n2418) );
  INV_X1 U1986 ( .A(\registers[4][6] ), .ZN(n2226) );
  INV_X1 U1987 ( .A(\registers[8][7] ), .ZN(n2289) );
  INV_X1 U1988 ( .A(\registers[14][7] ), .ZN(n2417) );
  INV_X1 U1989 ( .A(\registers[4][7] ), .ZN(n2225) );
  INV_X1 U1990 ( .A(\registers[8][8] ), .ZN(n2288) );
  INV_X1 U1991 ( .A(\registers[14][8] ), .ZN(n2416) );
  INV_X1 U1992 ( .A(\registers[4][8] ), .ZN(n2224) );
  INV_X1 U1993 ( .A(\registers[8][9] ), .ZN(n2287) );
  INV_X1 U1994 ( .A(\registers[14][9] ), .ZN(n2415) );
  INV_X1 U1995 ( .A(\registers[4][9] ), .ZN(n2223) );
  INV_X1 U1996 ( .A(\registers[8][10] ), .ZN(n2286) );
  INV_X1 U1997 ( .A(\registers[14][10] ), .ZN(n2414) );
  INV_X1 U1998 ( .A(\registers[4][10] ), .ZN(n2222) );
  INV_X1 U1999 ( .A(\registers[8][11] ), .ZN(n2285) );
  INV_X1 U2000 ( .A(\registers[14][11] ), .ZN(n2413) );
  INV_X1 U2001 ( .A(\registers[4][11] ), .ZN(n2221) );
  INV_X1 U2002 ( .A(\registers[8][12] ), .ZN(n2284) );
  INV_X1 U2003 ( .A(\registers[14][12] ), .ZN(n2412) );
  INV_X1 U2004 ( .A(\registers[4][12] ), .ZN(n2220) );
  INV_X1 U2005 ( .A(\registers[8][13] ), .ZN(n2283) );
  INV_X1 U2006 ( .A(\registers[14][13] ), .ZN(n2411) );
  INV_X1 U2007 ( .A(\registers[4][13] ), .ZN(n2219) );
  INV_X1 U2008 ( .A(\registers[8][14] ), .ZN(n2282) );
  INV_X1 U2009 ( .A(\registers[14][14] ), .ZN(n2410) );
  INV_X1 U2010 ( .A(\registers[4][14] ), .ZN(n2218) );
  INV_X1 U2011 ( .A(\registers[8][15] ), .ZN(n2281) );
  INV_X1 U2012 ( .A(\registers[14][15] ), .ZN(n2409) );
  INV_X1 U2013 ( .A(\registers[4][15] ), .ZN(n2217) );
  INV_X1 U2014 ( .A(\registers[8][16] ), .ZN(n2280) );
  INV_X1 U2015 ( .A(\registers[14][16] ), .ZN(n2408) );
  INV_X1 U2016 ( .A(\registers[4][16] ), .ZN(n2216) );
  INV_X1 U2017 ( .A(\registers[8][17] ), .ZN(n2279) );
  INV_X1 U2018 ( .A(\registers[14][17] ), .ZN(n2407) );
  INV_X1 U2019 ( .A(\registers[4][17] ), .ZN(n2215) );
  INV_X1 U2020 ( .A(\registers[8][18] ), .ZN(n2278) );
  INV_X1 U2021 ( .A(\registers[14][18] ), .ZN(n2406) );
  INV_X1 U2022 ( .A(\registers[4][18] ), .ZN(n2214) );
  INV_X1 U2023 ( .A(\registers[8][19] ), .ZN(n2277) );
  INV_X1 U2024 ( .A(\registers[14][19] ), .ZN(n2405) );
  INV_X1 U2025 ( .A(\registers[4][19] ), .ZN(n2213) );
  INV_X1 U2026 ( .A(\registers[8][20] ), .ZN(n2276) );
  INV_X1 U2027 ( .A(\registers[14][20] ), .ZN(n2404) );
  INV_X1 U2028 ( .A(\registers[4][20] ), .ZN(n2212) );
  INV_X1 U2029 ( .A(\registers[8][21] ), .ZN(n2275) );
  INV_X1 U2030 ( .A(\registers[14][21] ), .ZN(n2403) );
  INV_X1 U2031 ( .A(\registers[4][21] ), .ZN(n2211) );
  INV_X1 U2032 ( .A(\registers[8][22] ), .ZN(n2274) );
  INV_X1 U2033 ( .A(\registers[14][22] ), .ZN(n2402) );
  INV_X1 U2034 ( .A(\registers[4][22] ), .ZN(n2210) );
  INV_X1 U2035 ( .A(\registers[8][23] ), .ZN(n2273) );
  INV_X1 U2036 ( .A(\registers[14][23] ), .ZN(n2401) );
  INV_X1 U2037 ( .A(\registers[4][23] ), .ZN(n2209) );
  INV_X1 U2038 ( .A(\registers[8][24] ), .ZN(n2272) );
  INV_X1 U2039 ( .A(\registers[14][24] ), .ZN(n2400) );
  INV_X1 U2040 ( .A(\registers[4][24] ), .ZN(n2208) );
  INV_X1 U2041 ( .A(\registers[8][25] ), .ZN(n2271) );
  INV_X1 U2042 ( .A(\registers[14][25] ), .ZN(n2399) );
  INV_X1 U2043 ( .A(\registers[4][25] ), .ZN(n2207) );
  INV_X1 U2044 ( .A(\registers[8][26] ), .ZN(n2270) );
  INV_X1 U2045 ( .A(\registers[14][26] ), .ZN(n2398) );
  INV_X1 U2046 ( .A(\registers[4][26] ), .ZN(n2206) );
  INV_X1 U2047 ( .A(\registers[8][27] ), .ZN(n2269) );
  INV_X1 U2048 ( .A(\registers[14][27] ), .ZN(n2397) );
  INV_X1 U2049 ( .A(\registers[4][27] ), .ZN(n2205) );
  INV_X1 U2050 ( .A(\registers[8][28] ), .ZN(n2268) );
  INV_X1 U2051 ( .A(\registers[14][28] ), .ZN(n2396) );
  INV_X1 U2052 ( .A(\registers[4][28] ), .ZN(n2204) );
  INV_X1 U2053 ( .A(\registers[8][29] ), .ZN(n2267) );
  INV_X1 U2054 ( .A(\registers[14][29] ), .ZN(n2395) );
  INV_X1 U2055 ( .A(\registers[4][29] ), .ZN(n2203) );
  INV_X1 U2056 ( .A(\registers[8][30] ), .ZN(n2266) );
  INV_X1 U2057 ( .A(\registers[14][30] ), .ZN(n2394) );
  INV_X1 U2058 ( .A(\registers[4][30] ), .ZN(n2202) );
  INV_X1 U2059 ( .A(\registers[8][31] ), .ZN(n2265) );
  INV_X1 U2060 ( .A(\registers[14][31] ), .ZN(n2393) );
  INV_X1 U2061 ( .A(\registers[4][31] ), .ZN(n2201) );
  INV_X1 U2062 ( .A(\registers[18][0] ), .ZN(n2456) );
  INV_X1 U2063 ( .A(\registers[20][0] ), .ZN(n2520) );
  INV_X1 U2064 ( .A(\registers[26][0] ), .ZN(n2584) );
  INV_X1 U2065 ( .A(\registers[28][0] ), .ZN(n2648) );
  INV_X1 U2066 ( .A(\registers[7][0] ), .ZN(n2264) );
  INV_X1 U2067 ( .A(\registers[18][1] ), .ZN(n2455) );
  INV_X1 U2068 ( .A(\registers[20][1] ), .ZN(n2519) );
  INV_X1 U2069 ( .A(\registers[26][1] ), .ZN(n2583) );
  INV_X1 U2070 ( .A(\registers[28][1] ), .ZN(n2647) );
  INV_X1 U2071 ( .A(\registers[7][1] ), .ZN(n2263) );
  INV_X1 U2072 ( .A(\registers[18][2] ), .ZN(n2454) );
  INV_X1 U2073 ( .A(\registers[20][2] ), .ZN(n2518) );
  INV_X1 U2074 ( .A(\registers[26][2] ), .ZN(n2582) );
  INV_X1 U2075 ( .A(\registers[28][2] ), .ZN(n2646) );
  INV_X1 U2076 ( .A(\registers[7][2] ), .ZN(n2262) );
  INV_X1 U2077 ( .A(\registers[18][3] ), .ZN(n2453) );
  INV_X1 U2078 ( .A(\registers[20][3] ), .ZN(n2517) );
  INV_X1 U2079 ( .A(\registers[26][3] ), .ZN(n2581) );
  INV_X1 U2080 ( .A(\registers[28][3] ), .ZN(n2645) );
  INV_X1 U2081 ( .A(\registers[7][3] ), .ZN(n2261) );
  INV_X1 U2082 ( .A(\registers[18][4] ), .ZN(n2452) );
  INV_X1 U2083 ( .A(\registers[20][4] ), .ZN(n2516) );
  INV_X1 U2084 ( .A(\registers[26][4] ), .ZN(n2580) );
  INV_X1 U2085 ( .A(\registers[28][4] ), .ZN(n2644) );
  INV_X1 U2086 ( .A(\registers[7][4] ), .ZN(n2260) );
  INV_X1 U2087 ( .A(\registers[18][5] ), .ZN(n2451) );
  INV_X1 U2088 ( .A(\registers[20][5] ), .ZN(n2515) );
  INV_X1 U2089 ( .A(\registers[26][5] ), .ZN(n2579) );
  INV_X1 U2090 ( .A(\registers[28][5] ), .ZN(n2643) );
  INV_X1 U2091 ( .A(\registers[7][5] ), .ZN(n2259) );
  INV_X1 U2092 ( .A(\registers[18][6] ), .ZN(n2450) );
  INV_X1 U2093 ( .A(\registers[20][6] ), .ZN(n2514) );
  INV_X1 U2094 ( .A(\registers[26][6] ), .ZN(n2578) );
  INV_X1 U2095 ( .A(\registers[28][6] ), .ZN(n2642) );
  INV_X1 U2096 ( .A(\registers[7][6] ), .ZN(n2258) );
  INV_X1 U2097 ( .A(\registers[18][7] ), .ZN(n2449) );
  INV_X1 U2098 ( .A(\registers[20][7] ), .ZN(n2513) );
  INV_X1 U2099 ( .A(\registers[26][7] ), .ZN(n2577) );
  INV_X1 U2100 ( .A(\registers[28][7] ), .ZN(n2641) );
  INV_X1 U2101 ( .A(\registers[7][7] ), .ZN(n2257) );
  INV_X1 U2102 ( .A(\registers[18][8] ), .ZN(n2448) );
  INV_X1 U2103 ( .A(\registers[20][8] ), .ZN(n2512) );
  INV_X1 U2104 ( .A(\registers[26][8] ), .ZN(n2576) );
  INV_X1 U2105 ( .A(\registers[28][8] ), .ZN(n2640) );
  INV_X1 U2106 ( .A(\registers[7][8] ), .ZN(n2256) );
  INV_X1 U2107 ( .A(\registers[18][9] ), .ZN(n2447) );
  INV_X1 U2108 ( .A(\registers[20][9] ), .ZN(n2511) );
  INV_X1 U2109 ( .A(\registers[26][9] ), .ZN(n2575) );
  INV_X1 U2110 ( .A(\registers[28][9] ), .ZN(n2639) );
  INV_X1 U2111 ( .A(\registers[7][9] ), .ZN(n2255) );
  INV_X1 U2112 ( .A(\registers[18][10] ), .ZN(n2446) );
  INV_X1 U2113 ( .A(\registers[20][10] ), .ZN(n2510) );
  INV_X1 U2114 ( .A(\registers[26][10] ), .ZN(n2574) );
  INV_X1 U2115 ( .A(\registers[28][10] ), .ZN(n2638) );
  INV_X1 U2116 ( .A(\registers[7][10] ), .ZN(n2254) );
  INV_X1 U2117 ( .A(\registers[18][11] ), .ZN(n2445) );
  INV_X1 U2118 ( .A(\registers[20][11] ), .ZN(n2509) );
  INV_X1 U2119 ( .A(\registers[26][11] ), .ZN(n2573) );
  INV_X1 U2120 ( .A(\registers[28][11] ), .ZN(n2637) );
  INV_X1 U2121 ( .A(\registers[7][11] ), .ZN(n2253) );
  INV_X1 U2122 ( .A(\registers[18][12] ), .ZN(n2444) );
  INV_X1 U2123 ( .A(\registers[20][12] ), .ZN(n2508) );
  INV_X1 U2124 ( .A(\registers[26][12] ), .ZN(n2572) );
  INV_X1 U2125 ( .A(\registers[28][12] ), .ZN(n2636) );
  INV_X1 U2126 ( .A(\registers[7][12] ), .ZN(n2252) );
  INV_X1 U2127 ( .A(\registers[18][13] ), .ZN(n2443) );
  INV_X1 U2128 ( .A(\registers[20][13] ), .ZN(n2507) );
  INV_X1 U2129 ( .A(\registers[26][13] ), .ZN(n2571) );
  INV_X1 U2130 ( .A(\registers[28][13] ), .ZN(n2635) );
  INV_X1 U2131 ( .A(\registers[7][13] ), .ZN(n2251) );
  INV_X1 U2132 ( .A(\registers[18][14] ), .ZN(n2442) );
  INV_X1 U2133 ( .A(\registers[20][14] ), .ZN(n2506) );
  INV_X1 U2134 ( .A(\registers[26][14] ), .ZN(n2570) );
  INV_X1 U2135 ( .A(\registers[28][14] ), .ZN(n2634) );
  INV_X1 U2136 ( .A(\registers[7][14] ), .ZN(n2250) );
  INV_X1 U2137 ( .A(\registers[18][15] ), .ZN(n2441) );
  INV_X1 U2138 ( .A(\registers[20][15] ), .ZN(n2505) );
  INV_X1 U2139 ( .A(\registers[26][15] ), .ZN(n2569) );
  INV_X1 U2140 ( .A(\registers[28][15] ), .ZN(n2633) );
  INV_X1 U2141 ( .A(\registers[7][15] ), .ZN(n2249) );
  INV_X1 U2142 ( .A(\registers[18][16] ), .ZN(n2440) );
  INV_X1 U2143 ( .A(\registers[20][16] ), .ZN(n2504) );
  INV_X1 U2144 ( .A(\registers[26][16] ), .ZN(n2568) );
  INV_X1 U2145 ( .A(\registers[28][16] ), .ZN(n2632) );
  INV_X1 U2146 ( .A(\registers[7][16] ), .ZN(n2248) );
  INV_X1 U2147 ( .A(\registers[18][17] ), .ZN(n2439) );
  INV_X1 U2148 ( .A(\registers[20][17] ), .ZN(n2503) );
  INV_X1 U2149 ( .A(\registers[26][17] ), .ZN(n2567) );
  INV_X1 U2150 ( .A(\registers[28][17] ), .ZN(n2631) );
  INV_X1 U2151 ( .A(\registers[7][17] ), .ZN(n2247) );
  INV_X1 U2152 ( .A(\registers[18][18] ), .ZN(n2438) );
  INV_X1 U2153 ( .A(\registers[20][18] ), .ZN(n2502) );
  INV_X1 U2154 ( .A(\registers[26][18] ), .ZN(n2566) );
  INV_X1 U2155 ( .A(\registers[28][18] ), .ZN(n2630) );
  INV_X1 U2156 ( .A(\registers[7][18] ), .ZN(n2246) );
  INV_X1 U2157 ( .A(\registers[18][19] ), .ZN(n2437) );
  INV_X1 U2158 ( .A(\registers[20][19] ), .ZN(n2501) );
  INV_X1 U2159 ( .A(\registers[26][19] ), .ZN(n2565) );
  INV_X1 U2160 ( .A(\registers[28][19] ), .ZN(n2629) );
  INV_X1 U2161 ( .A(\registers[7][19] ), .ZN(n2245) );
  INV_X1 U2162 ( .A(\registers[18][20] ), .ZN(n2436) );
  INV_X1 U2163 ( .A(\registers[20][20] ), .ZN(n2500) );
  INV_X1 U2164 ( .A(\registers[26][20] ), .ZN(n2564) );
  INV_X1 U2165 ( .A(\registers[28][20] ), .ZN(n2628) );
  INV_X1 U2166 ( .A(\registers[7][20] ), .ZN(n2244) );
  INV_X1 U2167 ( .A(\registers[18][21] ), .ZN(n2435) );
  INV_X1 U2168 ( .A(\registers[20][21] ), .ZN(n2499) );
  INV_X1 U2169 ( .A(\registers[26][21] ), .ZN(n2563) );
  INV_X1 U2170 ( .A(\registers[28][21] ), .ZN(n2627) );
  INV_X1 U2171 ( .A(\registers[7][21] ), .ZN(n2243) );
  INV_X1 U2172 ( .A(\registers[18][22] ), .ZN(n2434) );
  INV_X1 U2173 ( .A(\registers[20][22] ), .ZN(n2498) );
  INV_X1 U2174 ( .A(\registers[26][22] ), .ZN(n2562) );
  INV_X1 U2175 ( .A(\registers[28][22] ), .ZN(n2626) );
  INV_X1 U2176 ( .A(\registers[7][22] ), .ZN(n2242) );
  INV_X1 U2177 ( .A(\registers[18][23] ), .ZN(n2433) );
  INV_X1 U2178 ( .A(\registers[20][23] ), .ZN(n2497) );
  INV_X1 U2179 ( .A(\registers[26][23] ), .ZN(n2561) );
  INV_X1 U2180 ( .A(\registers[28][23] ), .ZN(n2625) );
  INV_X1 U2181 ( .A(\registers[7][23] ), .ZN(n2241) );
  INV_X1 U2182 ( .A(\registers[18][24] ), .ZN(n2432) );
  INV_X1 U2183 ( .A(\registers[20][24] ), .ZN(n2496) );
  INV_X1 U2184 ( .A(\registers[26][24] ), .ZN(n2560) );
  INV_X1 U2185 ( .A(\registers[28][24] ), .ZN(n2624) );
  INV_X1 U2186 ( .A(\registers[7][24] ), .ZN(n2240) );
  INV_X1 U2187 ( .A(\registers[18][25] ), .ZN(n2431) );
  INV_X1 U2188 ( .A(\registers[20][25] ), .ZN(n2495) );
  INV_X1 U2189 ( .A(\registers[26][25] ), .ZN(n2559) );
  INV_X1 U2190 ( .A(\registers[28][25] ), .ZN(n2623) );
  INV_X1 U2191 ( .A(\registers[7][25] ), .ZN(n2239) );
  INV_X1 U2192 ( .A(\registers[18][26] ), .ZN(n2430) );
  INV_X1 U2193 ( .A(\registers[20][26] ), .ZN(n2494) );
  INV_X1 U2194 ( .A(\registers[26][26] ), .ZN(n2558) );
  INV_X1 U2195 ( .A(\registers[28][26] ), .ZN(n2622) );
  INV_X1 U2196 ( .A(\registers[7][26] ), .ZN(n2238) );
  INV_X1 U2197 ( .A(\registers[18][27] ), .ZN(n2429) );
  INV_X1 U2198 ( .A(\registers[20][27] ), .ZN(n2493) );
  INV_X1 U2199 ( .A(\registers[26][27] ), .ZN(n2557) );
  INV_X1 U2200 ( .A(\registers[28][27] ), .ZN(n2621) );
  INV_X1 U2201 ( .A(\registers[7][27] ), .ZN(n2237) );
  INV_X1 U2202 ( .A(\registers[18][28] ), .ZN(n2428) );
  INV_X1 U2203 ( .A(\registers[20][28] ), .ZN(n2492) );
  INV_X1 U2204 ( .A(\registers[26][28] ), .ZN(n2556) );
  INV_X1 U2205 ( .A(\registers[28][28] ), .ZN(n2620) );
  INV_X1 U2206 ( .A(\registers[7][28] ), .ZN(n2236) );
  INV_X1 U2207 ( .A(\registers[18][29] ), .ZN(n2427) );
  INV_X1 U2208 ( .A(\registers[20][29] ), .ZN(n2491) );
  INV_X1 U2209 ( .A(\registers[26][29] ), .ZN(n2555) );
  INV_X1 U2210 ( .A(\registers[28][29] ), .ZN(n2619) );
  INV_X1 U2211 ( .A(\registers[7][29] ), .ZN(n2235) );
  INV_X1 U2212 ( .A(\registers[18][30] ), .ZN(n2426) );
  INV_X1 U2213 ( .A(\registers[20][30] ), .ZN(n2490) );
  INV_X1 U2214 ( .A(\registers[26][30] ), .ZN(n2554) );
  INV_X1 U2215 ( .A(\registers[28][30] ), .ZN(n2618) );
  INV_X1 U2216 ( .A(\registers[7][30] ), .ZN(n2234) );
  INV_X1 U2217 ( .A(\registers[18][31] ), .ZN(n2425) );
  INV_X1 U2218 ( .A(\registers[20][31] ), .ZN(n2489) );
  INV_X1 U2219 ( .A(\registers[26][31] ), .ZN(n2553) );
  INV_X1 U2220 ( .A(\registers[28][31] ), .ZN(n2617) );
  INV_X1 U2221 ( .A(\registers[7][31] ), .ZN(n2233) );
  INV_X1 U2222 ( .A(add_wr[4]), .ZN(n2164) );
  INV_X1 U2223 ( .A(add_wr[3]), .ZN(n2165) );
  AND2_X1 U2224 ( .A1(wr), .A2(n2689), .ZN(n535) );
  INV_X1 U2225 ( .A(enable), .ZN(n2689) );
  CLKBUF_X1 U2226 ( .A(N371), .Z(n1962) );
  CLKBUF_X1 U2227 ( .A(N371), .Z(n1963) );
  CLKBUF_X1 U2228 ( .A(N371), .Z(n1964) );
  CLKBUF_X1 U2229 ( .A(N371), .Z(n1965) );
  CLKBUF_X1 U2230 ( .A(N371), .Z(n1966) );
  CLKBUF_X1 U2231 ( .A(N371), .Z(n1967) );
endmodule


module sign_extension_sign_init16_sign_ext32 ( data_in, data_out );
  input [15:0] data_in;
  output [31:0] data_out;
  wire   data_out_31;
  assign data_out[31] = data_out_31;
  assign data_out[30] = data_out_31;
  assign data_out[29] = data_out_31;
  assign data_out[28] = data_out_31;
  assign data_out[27] = data_out_31;
  assign data_out[26] = data_out_31;
  assign data_out[25] = data_out_31;
  assign data_out[24] = data_out_31;
  assign data_out[23] = data_out_31;
  assign data_out[22] = data_out_31;
  assign data_out[21] = data_out_31;
  assign data_out[20] = data_out_31;
  assign data_out[19] = data_out_31;
  assign data_out[18] = data_out_31;
  assign data_out[17] = data_out_31;
  assign data_out[16] = data_out_31;
  assign data_out[15] = data_out_31;
  assign data_out_31 = data_in[15];
  assign data_out[14] = data_in[14];
  assign data_out[13] = data_in[13];
  assign data_out[12] = data_in[12];
  assign data_out[11] = data_in[11];
  assign data_out[10] = data_in[10];
  assign data_out[9] = data_in[9];
  assign data_out[8] = data_in[8];
  assign data_out[7] = data_in[7];
  assign data_out[6] = data_in[6];
  assign data_out[5] = data_in[5];
  assign data_out[4] = data_in[4];
  assign data_out[3] = data_in[3];
  assign data_out[2] = data_in[2];
  assign data_out[1] = data_in[1];
  assign data_out[0] = data_in[0];

endmodule


module REG_GEN_NBIT32_16 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n52), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n52), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n52), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n52), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n52), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n52), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n52), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n52), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n51), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n51), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n51), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n51), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n51), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n51), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n51), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n50), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n50), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n50), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n50), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n50), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n50), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n50), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n50), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n50), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n50), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n50), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n50), .Q(Q[0]), .QN(n97) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n36), .Z(n42) );
  BUF_X1 U10 ( .A(n37), .Z(n44) );
  BUF_X1 U11 ( .A(n37), .Z(n45) );
  BUF_X1 U12 ( .A(n37), .Z(n46) );
  BUF_X1 U13 ( .A(n38), .Z(n47) );
  BUF_X1 U14 ( .A(n38), .Z(n48) );
  BUF_X1 U15 ( .A(n36), .Z(n41) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n36) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n37) );
  OAI22_X1 U19 ( .A1(n97), .A2(n39), .B1(n42), .B2(n57), .ZN(n35) );
  INV_X1 U20 ( .A(D[0]), .ZN(n57) );
  OAI22_X1 U21 ( .A1(n96), .A2(n40), .B1(n42), .B2(n56), .ZN(n34) );
  INV_X1 U22 ( .A(D[1]), .ZN(n56) );
  OAI22_X1 U23 ( .A1(n71), .A2(n40), .B1(n41), .B2(n111), .ZN(n9) );
  INV_X1 U24 ( .A(D[26]), .ZN(n111) );
  OAI22_X1 U25 ( .A1(n70), .A2(n39), .B1(n41), .B2(n112), .ZN(n8) );
  INV_X1 U26 ( .A(D[27]), .ZN(n112) );
  OAI22_X1 U27 ( .A1(n69), .A2(n40), .B1(n41), .B2(n113), .ZN(n7) );
  INV_X1 U28 ( .A(D[28]), .ZN(n113) );
  OAI22_X1 U29 ( .A1(n68), .A2(n39), .B1(n41), .B2(n114), .ZN(n6) );
  INV_X1 U30 ( .A(D[29]), .ZN(n114) );
  OAI22_X1 U31 ( .A1(n67), .A2(n40), .B1(n42), .B2(n115), .ZN(n5) );
  INV_X1 U32 ( .A(D[30]), .ZN(n115) );
  OAI22_X1 U33 ( .A1(n66), .A2(n39), .B1(n42), .B2(n116), .ZN(n4) );
  INV_X1 U34 ( .A(D[31]), .ZN(n116) );
  OAI22_X1 U35 ( .A1(n93), .A2(n40), .B1(n43), .B2(n53), .ZN(n31) );
  INV_X1 U36 ( .A(D[4]), .ZN(n53) );
  OAI22_X1 U37 ( .A1(n95), .A2(n40), .B1(n43), .B2(n55), .ZN(n33) );
  INV_X1 U38 ( .A(D[2]), .ZN(n55) );
  OAI22_X1 U39 ( .A1(n94), .A2(n40), .B1(n43), .B2(n54), .ZN(n32) );
  INV_X1 U40 ( .A(D[3]), .ZN(n54) );
  OAI22_X1 U41 ( .A1(n92), .A2(n40), .B1(n43), .B2(n58), .ZN(n30) );
  INV_X1 U42 ( .A(D[5]), .ZN(n58) );
  OAI22_X1 U43 ( .A1(n91), .A2(n40), .B1(n44), .B2(n59), .ZN(n29) );
  INV_X1 U44 ( .A(D[6]), .ZN(n59) );
  OAI22_X1 U45 ( .A1(n90), .A2(n40), .B1(n44), .B2(n60), .ZN(n28) );
  INV_X1 U46 ( .A(D[7]), .ZN(n60) );
  OAI22_X1 U47 ( .A1(n89), .A2(n40), .B1(n44), .B2(n61), .ZN(n27) );
  INV_X1 U48 ( .A(D[8]), .ZN(n61) );
  OAI22_X1 U49 ( .A1(n88), .A2(n40), .B1(n44), .B2(n62), .ZN(n26) );
  INV_X1 U50 ( .A(D[9]), .ZN(n62) );
  OAI22_X1 U51 ( .A1(n87), .A2(n40), .B1(n45), .B2(n63), .ZN(n25) );
  INV_X1 U52 ( .A(D[10]), .ZN(n63) );
  OAI22_X1 U53 ( .A1(n86), .A2(n40), .B1(n45), .B2(n64), .ZN(n24) );
  INV_X1 U54 ( .A(D[11]), .ZN(n64) );
  OAI22_X1 U55 ( .A1(n85), .A2(n40), .B1(n45), .B2(n65), .ZN(n23) );
  INV_X1 U56 ( .A(D[12]), .ZN(n65) );
  OAI22_X1 U57 ( .A1(n84), .A2(n40), .B1(n45), .B2(n98), .ZN(n22) );
  INV_X1 U58 ( .A(D[13]), .ZN(n98) );
  OAI22_X1 U59 ( .A1(n83), .A2(n39), .B1(n46), .B2(n99), .ZN(n21) );
  INV_X1 U60 ( .A(D[14]), .ZN(n99) );
  OAI22_X1 U61 ( .A1(n82), .A2(n39), .B1(n46), .B2(n100), .ZN(n20) );
  INV_X1 U62 ( .A(D[15]), .ZN(n100) );
  OAI22_X1 U63 ( .A1(n81), .A2(n39), .B1(n46), .B2(n101), .ZN(n19) );
  INV_X1 U64 ( .A(D[16]), .ZN(n101) );
  OAI22_X1 U65 ( .A1(n80), .A2(n39), .B1(n46), .B2(n102), .ZN(n18) );
  INV_X1 U66 ( .A(D[17]), .ZN(n102) );
  OAI22_X1 U67 ( .A1(n79), .A2(n39), .B1(n47), .B2(n103), .ZN(n17) );
  INV_X1 U68 ( .A(D[18]), .ZN(n103) );
  OAI22_X1 U69 ( .A1(n78), .A2(n39), .B1(n47), .B2(n104), .ZN(n16) );
  INV_X1 U70 ( .A(D[19]), .ZN(n104) );
  OAI22_X1 U71 ( .A1(n77), .A2(n39), .B1(n47), .B2(n105), .ZN(n15) );
  INV_X1 U72 ( .A(D[20]), .ZN(n105) );
  OAI22_X1 U73 ( .A1(n76), .A2(n39), .B1(n47), .B2(n106), .ZN(n14) );
  INV_X1 U74 ( .A(D[21]), .ZN(n106) );
  OAI22_X1 U75 ( .A1(n75), .A2(n39), .B1(n48), .B2(n107), .ZN(n13) );
  INV_X1 U76 ( .A(D[22]), .ZN(n107) );
  OAI22_X1 U77 ( .A1(n74), .A2(n39), .B1(n48), .B2(n108), .ZN(n12) );
  INV_X1 U78 ( .A(D[23]), .ZN(n108) );
  OAI22_X1 U79 ( .A1(n73), .A2(n39), .B1(n48), .B2(n109), .ZN(n11) );
  INV_X1 U80 ( .A(D[24]), .ZN(n109) );
  OAI22_X1 U81 ( .A1(n72), .A2(n39), .B1(n48), .B2(n110), .ZN(n10) );
  INV_X1 U82 ( .A(D[25]), .ZN(n110) );
endmodule


module REG_GEN_NBIT32_15 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n53), .Q(Q[31]), .QN(n149) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n53), .Q(Q[30]), .QN(n148) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n53), .Q(Q[29]), .QN(n147) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n53), .Q(Q[28]), .QN(n146) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n53), .Q(Q[27]), .QN(n145) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n53), .Q(Q[26]), .QN(n144) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n53), .Q(Q[25]), .QN(n143) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n53), .Q(Q[24]), .QN(n142) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n52), .Q(Q[23]), .QN(n141) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n52), .Q(Q[22]), .QN(n140) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n52), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n52), .Q(Q[20]), .QN(n138) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n52), .Q(Q[19]), .QN(n137) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n52), .Q(Q[18]), .QN(n136) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n52), .Q(Q[17]), .QN(n135) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n52), .Q(Q[16]), .QN(n134) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n52), .Q(Q[15]), .QN(n133) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n52), .Q(Q[14]), .QN(n132) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n52), .Q(Q[13]), .QN(n131) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n52), .Q(Q[12]), .QN(n130) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n51), .Q(Q[11]), .QN(n129) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n51), .Q(Q[10]), .QN(n128) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n51), .Q(Q[9]), .QN(n127) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n51), .Q(Q[8]), .QN(n126) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n51), .Q(Q[7]), .QN(n125) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n51), .Q(Q[6]), .QN(n124) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n51), .Q(Q[5]), .QN(n123) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n51), .Q(Q[4]), .QN(n122) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n51), .Q(Q[3]), .QN(n121) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n51), .Q(Q[2]), .QN(n120) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n51), .Q(Q[1]), .QN(n119) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n51), .Q(Q[0]), .QN(n118) );
  INV_X1 U2 ( .A(n50), .ZN(n40) );
  INV_X1 U3 ( .A(n50), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n53) );
  BUF_X1 U7 ( .A(n38), .Z(n50) );
  BUF_X1 U8 ( .A(n36), .Z(n44) );
  BUF_X1 U9 ( .A(n36), .Z(n43) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n37), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n38), .Z(n49) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n36) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n37) );
  OAI22_X1 U19 ( .A1(n118), .A2(n41), .B1(n43), .B2(n58), .ZN(n35) );
  INV_X1 U20 ( .A(D[0]), .ZN(n58) );
  OAI22_X1 U21 ( .A1(n119), .A2(n41), .B1(n43), .B2(n57), .ZN(n34) );
  INV_X1 U22 ( .A(D[1]), .ZN(n57) );
  OAI22_X1 U23 ( .A1(n144), .A2(n41), .B1(n42), .B2(n112), .ZN(n9) );
  INV_X1 U24 ( .A(D[26]), .ZN(n112) );
  OAI22_X1 U25 ( .A1(n145), .A2(n41), .B1(n42), .B2(n113), .ZN(n8) );
  INV_X1 U26 ( .A(D[27]), .ZN(n113) );
  OAI22_X1 U27 ( .A1(n146), .A2(n41), .B1(n42), .B2(n114), .ZN(n7) );
  INV_X1 U28 ( .A(D[28]), .ZN(n114) );
  OAI22_X1 U29 ( .A1(n147), .A2(n41), .B1(n42), .B2(n115), .ZN(n6) );
  INV_X1 U30 ( .A(D[29]), .ZN(n115) );
  OAI22_X1 U31 ( .A1(n148), .A2(n41), .B1(n43), .B2(n116), .ZN(n5) );
  INV_X1 U32 ( .A(D[30]), .ZN(n116) );
  OAI22_X1 U33 ( .A1(n149), .A2(n41), .B1(n43), .B2(n117), .ZN(n4) );
  INV_X1 U34 ( .A(D[31]), .ZN(n117) );
  OAI22_X1 U35 ( .A1(n120), .A2(n40), .B1(n44), .B2(n56), .ZN(n33) );
  INV_X1 U36 ( .A(D[2]), .ZN(n56) );
  OAI22_X1 U37 ( .A1(n121), .A2(n40), .B1(n44), .B2(n55), .ZN(n32) );
  INV_X1 U38 ( .A(D[3]), .ZN(n55) );
  OAI22_X1 U39 ( .A1(n122), .A2(n40), .B1(n44), .B2(n54), .ZN(n31) );
  INV_X1 U40 ( .A(D[4]), .ZN(n54) );
  OAI22_X1 U41 ( .A1(n123), .A2(n40), .B1(n44), .B2(n59), .ZN(n30) );
  INV_X1 U42 ( .A(D[5]), .ZN(n59) );
  OAI22_X1 U43 ( .A1(n124), .A2(n40), .B1(n45), .B2(n60), .ZN(n29) );
  INV_X1 U44 ( .A(D[6]), .ZN(n60) );
  OAI22_X1 U45 ( .A1(n125), .A2(n40), .B1(n45), .B2(n61), .ZN(n28) );
  INV_X1 U46 ( .A(D[7]), .ZN(n61) );
  OAI22_X1 U47 ( .A1(n126), .A2(n40), .B1(n45), .B2(n62), .ZN(n27) );
  INV_X1 U48 ( .A(D[8]), .ZN(n62) );
  OAI22_X1 U49 ( .A1(n127), .A2(n40), .B1(n45), .B2(n63), .ZN(n26) );
  INV_X1 U50 ( .A(D[9]), .ZN(n63) );
  OAI22_X1 U51 ( .A1(n128), .A2(n40), .B1(n46), .B2(n64), .ZN(n25) );
  INV_X1 U52 ( .A(D[10]), .ZN(n64) );
  OAI22_X1 U53 ( .A1(n129), .A2(n40), .B1(n46), .B2(n65), .ZN(n24) );
  INV_X1 U54 ( .A(D[11]), .ZN(n65) );
  OAI22_X1 U55 ( .A1(n130), .A2(n40), .B1(n46), .B2(n98), .ZN(n23) );
  INV_X1 U56 ( .A(D[12]), .ZN(n98) );
  OAI22_X1 U57 ( .A1(n131), .A2(n40), .B1(n46), .B2(n99), .ZN(n22) );
  INV_X1 U58 ( .A(D[13]), .ZN(n99) );
  OAI22_X1 U59 ( .A1(n132), .A2(n39), .B1(n47), .B2(n100), .ZN(n21) );
  INV_X1 U60 ( .A(D[14]), .ZN(n100) );
  OAI22_X1 U61 ( .A1(n133), .A2(n39), .B1(n47), .B2(n101), .ZN(n20) );
  INV_X1 U62 ( .A(D[15]), .ZN(n101) );
  OAI22_X1 U63 ( .A1(n134), .A2(n39), .B1(n47), .B2(n102), .ZN(n19) );
  INV_X1 U64 ( .A(D[16]), .ZN(n102) );
  OAI22_X1 U65 ( .A1(n135), .A2(n39), .B1(n47), .B2(n103), .ZN(n18) );
  INV_X1 U66 ( .A(D[17]), .ZN(n103) );
  OAI22_X1 U67 ( .A1(n136), .A2(n39), .B1(n48), .B2(n104), .ZN(n17) );
  INV_X1 U68 ( .A(D[18]), .ZN(n104) );
  OAI22_X1 U69 ( .A1(n137), .A2(n39), .B1(n48), .B2(n105), .ZN(n16) );
  INV_X1 U70 ( .A(D[19]), .ZN(n105) );
  OAI22_X1 U71 ( .A1(n138), .A2(n39), .B1(n48), .B2(n106), .ZN(n15) );
  INV_X1 U72 ( .A(D[20]), .ZN(n106) );
  OAI22_X1 U73 ( .A1(n139), .A2(n39), .B1(n48), .B2(n107), .ZN(n14) );
  INV_X1 U74 ( .A(D[21]), .ZN(n107) );
  OAI22_X1 U75 ( .A1(n140), .A2(n39), .B1(n49), .B2(n108), .ZN(n13) );
  INV_X1 U76 ( .A(D[22]), .ZN(n108) );
  OAI22_X1 U77 ( .A1(n141), .A2(n39), .B1(n49), .B2(n109), .ZN(n12) );
  INV_X1 U78 ( .A(D[23]), .ZN(n109) );
  OAI22_X1 U79 ( .A1(n142), .A2(n39), .B1(n49), .B2(n110), .ZN(n11) );
  INV_X1 U80 ( .A(D[24]), .ZN(n110) );
  OAI22_X1 U81 ( .A1(n143), .A2(n39), .B1(n49), .B2(n111), .ZN(n10) );
  INV_X1 U82 ( .A(D[25]), .ZN(n111) );
  INV_X1 U83 ( .A(n50), .ZN(n41) );
endmodule


module REG_GEN_NBIT32_14 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n51), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n51), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n51), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n51), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n51), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n51), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n51), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n52), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n52), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n52), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n52), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n52), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n52), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n52), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n51), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n51), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n50), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n50), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n50), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n50), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n50), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n50), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n50), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n50), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n50), .Q(Q[0]), .QN(n97) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n51), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n50), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n51), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n52), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n50), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n50), .Q(Q[2]), .QN(n95) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n44) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n71), .A2(n40), .B1(n41), .B2(n64), .ZN(n9) );
  INV_X1 U20 ( .A(D[26]), .ZN(n64) );
  OAI22_X1 U21 ( .A1(n68), .A2(n39), .B1(n41), .B2(n99), .ZN(n6) );
  INV_X1 U22 ( .A(D[29]), .ZN(n99) );
  OAI22_X1 U23 ( .A1(n70), .A2(n40), .B1(n41), .B2(n65), .ZN(n8) );
  INV_X1 U24 ( .A(D[27]), .ZN(n65) );
  OAI22_X1 U25 ( .A1(n69), .A2(n39), .B1(n41), .B2(n98), .ZN(n7) );
  INV_X1 U26 ( .A(D[28]), .ZN(n98) );
  OAI22_X1 U27 ( .A1(n67), .A2(n40), .B1(n42), .B2(n100), .ZN(n5) );
  INV_X1 U28 ( .A(D[30]), .ZN(n100) );
  OAI22_X1 U29 ( .A1(n66), .A2(n39), .B1(n42), .B2(n101), .ZN(n4) );
  INV_X1 U30 ( .A(D[31]), .ZN(n101) );
  OAI22_X1 U31 ( .A1(n96), .A2(n40), .B1(n42), .B2(n115), .ZN(n34) );
  INV_X1 U32 ( .A(D[1]), .ZN(n115) );
  OAI22_X1 U33 ( .A1(n97), .A2(n39), .B1(n42), .B2(n116), .ZN(n35) );
  INV_X1 U34 ( .A(D[0]), .ZN(n116) );
  OAI22_X1 U35 ( .A1(n82), .A2(n39), .B1(n46), .B2(n53), .ZN(n20) );
  INV_X1 U36 ( .A(D[15]), .ZN(n53) );
  OAI22_X1 U37 ( .A1(n81), .A2(n39), .B1(n46), .B2(n54), .ZN(n19) );
  INV_X1 U38 ( .A(D[16]), .ZN(n54) );
  OAI22_X1 U39 ( .A1(n80), .A2(n39), .B1(n46), .B2(n55), .ZN(n18) );
  INV_X1 U40 ( .A(D[17]), .ZN(n55) );
  OAI22_X1 U41 ( .A1(n79), .A2(n39), .B1(n47), .B2(n56), .ZN(n17) );
  INV_X1 U42 ( .A(D[18]), .ZN(n56) );
  OAI22_X1 U43 ( .A1(n78), .A2(n39), .B1(n47), .B2(n57), .ZN(n16) );
  INV_X1 U44 ( .A(D[19]), .ZN(n57) );
  OAI22_X1 U45 ( .A1(n77), .A2(n39), .B1(n47), .B2(n58), .ZN(n15) );
  INV_X1 U46 ( .A(D[20]), .ZN(n58) );
  OAI22_X1 U47 ( .A1(n76), .A2(n39), .B1(n47), .B2(n59), .ZN(n14) );
  INV_X1 U48 ( .A(D[21]), .ZN(n59) );
  OAI22_X1 U49 ( .A1(n75), .A2(n39), .B1(n48), .B2(n60), .ZN(n13) );
  INV_X1 U50 ( .A(D[22]), .ZN(n60) );
  OAI22_X1 U51 ( .A1(n74), .A2(n39), .B1(n48), .B2(n61), .ZN(n12) );
  INV_X1 U52 ( .A(D[23]), .ZN(n61) );
  OAI22_X1 U53 ( .A1(n73), .A2(n39), .B1(n48), .B2(n62), .ZN(n11) );
  INV_X1 U54 ( .A(D[24]), .ZN(n62) );
  OAI22_X1 U55 ( .A1(n72), .A2(n39), .B1(n48), .B2(n63), .ZN(n10) );
  INV_X1 U56 ( .A(D[25]), .ZN(n63) );
  OAI22_X1 U57 ( .A1(n91), .A2(n40), .B1(n44), .B2(n110), .ZN(n29) );
  INV_X1 U58 ( .A(D[6]), .ZN(n110) );
  OAI22_X1 U59 ( .A1(n90), .A2(n40), .B1(n44), .B2(n109), .ZN(n28) );
  INV_X1 U60 ( .A(D[7]), .ZN(n109) );
  OAI22_X1 U61 ( .A1(n89), .A2(n40), .B1(n44), .B2(n108), .ZN(n27) );
  INV_X1 U62 ( .A(D[8]), .ZN(n108) );
  OAI22_X1 U63 ( .A1(n88), .A2(n40), .B1(n44), .B2(n107), .ZN(n26) );
  INV_X1 U64 ( .A(D[9]), .ZN(n107) );
  OAI22_X1 U65 ( .A1(n87), .A2(n40), .B1(n45), .B2(n106), .ZN(n25) );
  INV_X1 U66 ( .A(D[10]), .ZN(n106) );
  OAI22_X1 U67 ( .A1(n86), .A2(n40), .B1(n45), .B2(n105), .ZN(n24) );
  INV_X1 U68 ( .A(D[11]), .ZN(n105) );
  OAI22_X1 U69 ( .A1(n85), .A2(n40), .B1(n45), .B2(n104), .ZN(n23) );
  INV_X1 U70 ( .A(D[12]), .ZN(n104) );
  OAI22_X1 U71 ( .A1(n84), .A2(n40), .B1(n45), .B2(n103), .ZN(n22) );
  INV_X1 U72 ( .A(D[13]), .ZN(n103) );
  OAI22_X1 U73 ( .A1(n83), .A2(n39), .B1(n46), .B2(n102), .ZN(n21) );
  INV_X1 U74 ( .A(D[14]), .ZN(n102) );
  OAI22_X1 U75 ( .A1(n94), .A2(n40), .B1(n43), .B2(n113), .ZN(n32) );
  INV_X1 U76 ( .A(D[3]), .ZN(n113) );
  OAI22_X1 U77 ( .A1(n93), .A2(n40), .B1(n43), .B2(n112), .ZN(n31) );
  INV_X1 U78 ( .A(D[4]), .ZN(n112) );
  OAI22_X1 U79 ( .A1(n95), .A2(n40), .B1(n43), .B2(n114), .ZN(n33) );
  INV_X1 U80 ( .A(D[2]), .ZN(n114) );
  OAI22_X1 U81 ( .A1(n92), .A2(n40), .B1(n43), .B2(n111), .ZN(n30) );
  INV_X1 U82 ( .A(D[5]), .ZN(n111) );
endmodule


module REG_GEN_NBIT32_13 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n53), .Q(Q[31]), .QN(n149) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n53), .Q(Q[30]), .QN(n148) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n53), .Q(Q[29]), .QN(n147) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n53), .Q(Q[28]), .QN(n146) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n53), .Q(Q[27]), .QN(n145) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n53), .Q(Q[26]), .QN(n144) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n53), .Q(Q[25]), .QN(n143) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n53), .Q(Q[24]), .QN(n142) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n52), .Q(Q[23]), .QN(n141) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n52), .Q(Q[22]), .QN(n140) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n52), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n52), .Q(Q[20]), .QN(n138) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n52), .Q(Q[19]), .QN(n137) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n52), .Q(Q[18]), .QN(n136) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n52), .Q(Q[17]), .QN(n135) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n52), .Q(Q[16]), .QN(n134) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n52), .Q(Q[15]), .QN(n133) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n52), .Q(Q[14]), .QN(n132) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n52), .Q(Q[13]), .QN(n131) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n52), .Q(Q[12]), .QN(n130) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n51), .Q(Q[11]), .QN(n129) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n51), .Q(Q[10]), .QN(n128) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n51), .Q(Q[9]), .QN(n127) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n51), .Q(Q[8]), .QN(n126) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n51), .Q(Q[7]), .QN(n125) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n51), .Q(Q[6]), .QN(n124) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n51), .Q(Q[5]), .QN(n123) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n51), .Q(Q[4]), .QN(n122) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n51), .Q(Q[3]), .QN(n121) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n51), .Q(Q[2]), .QN(n120) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n51), .Q(Q[1]), .QN(n119) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n51), .Q(Q[0]), .QN(n118) );
  INV_X1 U2 ( .A(n50), .ZN(n40) );
  INV_X1 U3 ( .A(n50), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n53) );
  BUF_X1 U7 ( .A(n38), .Z(n50) );
  BUF_X1 U8 ( .A(n36), .Z(n44) );
  BUF_X1 U9 ( .A(n37), .Z(n45) );
  BUF_X1 U10 ( .A(n37), .Z(n46) );
  BUF_X1 U11 ( .A(n37), .Z(n47) );
  BUF_X1 U12 ( .A(n38), .Z(n48) );
  BUF_X1 U13 ( .A(n38), .Z(n49) );
  BUF_X1 U14 ( .A(n36), .Z(n42) );
  BUF_X1 U15 ( .A(n36), .Z(n43) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n144), .A2(n41), .B1(n42), .B2(n55), .ZN(n9) );
  INV_X1 U20 ( .A(D[26]), .ZN(n55) );
  OAI22_X1 U21 ( .A1(n145), .A2(n41), .B1(n42), .B2(n56), .ZN(n8) );
  INV_X1 U22 ( .A(D[27]), .ZN(n56) );
  OAI22_X1 U23 ( .A1(n146), .A2(n41), .B1(n42), .B2(n57), .ZN(n7) );
  INV_X1 U24 ( .A(D[28]), .ZN(n57) );
  OAI22_X1 U25 ( .A1(n147), .A2(n41), .B1(n42), .B2(n58), .ZN(n6) );
  INV_X1 U26 ( .A(D[29]), .ZN(n58) );
  OAI22_X1 U27 ( .A1(n148), .A2(n41), .B1(n43), .B2(n59), .ZN(n5) );
  INV_X1 U28 ( .A(D[30]), .ZN(n59) );
  OAI22_X1 U29 ( .A1(n149), .A2(n41), .B1(n43), .B2(n60), .ZN(n4) );
  INV_X1 U30 ( .A(D[31]), .ZN(n60) );
  OAI22_X1 U31 ( .A1(n119), .A2(n41), .B1(n43), .B2(n116), .ZN(n34) );
  INV_X1 U32 ( .A(D[1]), .ZN(n116) );
  OAI22_X1 U33 ( .A1(n118), .A2(n41), .B1(n43), .B2(n117), .ZN(n35) );
  INV_X1 U34 ( .A(D[0]), .ZN(n117) );
  OAI22_X1 U35 ( .A1(n133), .A2(n39), .B1(n47), .B2(n102), .ZN(n20) );
  INV_X1 U36 ( .A(D[15]), .ZN(n102) );
  OAI22_X1 U37 ( .A1(n143), .A2(n39), .B1(n49), .B2(n54), .ZN(n10) );
  INV_X1 U38 ( .A(D[25]), .ZN(n54) );
  OAI22_X1 U39 ( .A1(n122), .A2(n40), .B1(n44), .B2(n113), .ZN(n31) );
  INV_X1 U40 ( .A(D[4]), .ZN(n113) );
  OAI22_X1 U41 ( .A1(n126), .A2(n40), .B1(n45), .B2(n109), .ZN(n27) );
  INV_X1 U42 ( .A(D[8]), .ZN(n109) );
  OAI22_X1 U43 ( .A1(n127), .A2(n40), .B1(n45), .B2(n108), .ZN(n26) );
  INV_X1 U44 ( .A(D[9]), .ZN(n108) );
  OAI22_X1 U45 ( .A1(n128), .A2(n40), .B1(n46), .B2(n107), .ZN(n25) );
  INV_X1 U46 ( .A(D[10]), .ZN(n107) );
  OAI22_X1 U47 ( .A1(n129), .A2(n40), .B1(n46), .B2(n106), .ZN(n24) );
  INV_X1 U48 ( .A(D[11]), .ZN(n106) );
  OAI22_X1 U49 ( .A1(n130), .A2(n40), .B1(n46), .B2(n105), .ZN(n23) );
  INV_X1 U50 ( .A(D[12]), .ZN(n105) );
  OAI22_X1 U51 ( .A1(n131), .A2(n40), .B1(n46), .B2(n104), .ZN(n22) );
  INV_X1 U52 ( .A(D[13]), .ZN(n104) );
  OAI22_X1 U53 ( .A1(n132), .A2(n39), .B1(n47), .B2(n103), .ZN(n21) );
  INV_X1 U54 ( .A(D[14]), .ZN(n103) );
  OAI22_X1 U55 ( .A1(n120), .A2(n40), .B1(n44), .B2(n115), .ZN(n33) );
  INV_X1 U56 ( .A(D[2]), .ZN(n115) );
  OAI22_X1 U57 ( .A1(n121), .A2(n40), .B1(n44), .B2(n114), .ZN(n32) );
  INV_X1 U58 ( .A(D[3]), .ZN(n114) );
  OAI22_X1 U59 ( .A1(n123), .A2(n40), .B1(n44), .B2(n112), .ZN(n30) );
  INV_X1 U60 ( .A(D[5]), .ZN(n112) );
  OAI22_X1 U61 ( .A1(n124), .A2(n40), .B1(n45), .B2(n111), .ZN(n29) );
  INV_X1 U62 ( .A(D[6]), .ZN(n111) );
  OAI22_X1 U63 ( .A1(n125), .A2(n40), .B1(n45), .B2(n110), .ZN(n28) );
  INV_X1 U64 ( .A(D[7]), .ZN(n110) );
  OAI22_X1 U65 ( .A1(n134), .A2(n39), .B1(n47), .B2(n101), .ZN(n19) );
  INV_X1 U66 ( .A(D[16]), .ZN(n101) );
  OAI22_X1 U67 ( .A1(n135), .A2(n39), .B1(n47), .B2(n100), .ZN(n18) );
  INV_X1 U68 ( .A(D[17]), .ZN(n100) );
  OAI22_X1 U69 ( .A1(n136), .A2(n39), .B1(n48), .B2(n99), .ZN(n17) );
  INV_X1 U70 ( .A(D[18]), .ZN(n99) );
  OAI22_X1 U71 ( .A1(n137), .A2(n39), .B1(n48), .B2(n98), .ZN(n16) );
  INV_X1 U72 ( .A(D[19]), .ZN(n98) );
  OAI22_X1 U73 ( .A1(n139), .A2(n39), .B1(n48), .B2(n64), .ZN(n14) );
  INV_X1 U74 ( .A(D[21]), .ZN(n64) );
  OAI22_X1 U75 ( .A1(n140), .A2(n39), .B1(n49), .B2(n63), .ZN(n13) );
  INV_X1 U76 ( .A(D[22]), .ZN(n63) );
  OAI22_X1 U77 ( .A1(n141), .A2(n39), .B1(n49), .B2(n62), .ZN(n12) );
  INV_X1 U78 ( .A(D[23]), .ZN(n62) );
  OAI22_X1 U79 ( .A1(n142), .A2(n39), .B1(n49), .B2(n61), .ZN(n11) );
  INV_X1 U80 ( .A(D[24]), .ZN(n61) );
  OAI22_X1 U81 ( .A1(n138), .A2(n39), .B1(n48), .B2(n65), .ZN(n15) );
  INV_X1 U82 ( .A(D[20]), .ZN(n65) );
  INV_X1 U83 ( .A(n50), .ZN(n41) );
endmodule


module REG_GEN_NBIT32_12 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116;

  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n52), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n52), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n52), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n52), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n52), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n51), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n51), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n51), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n51), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n50), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n51), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n51), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n50), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n51), .Q(Q[0]), .QN(n97) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n50), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n50), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n52), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n52), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n50), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n50), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n51), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n52), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n50), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n50), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n50), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n51), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n50), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n50), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n50), .Q(Q[12]), .QN(n85) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n37), .Z(n44) );
  BUF_X1 U9 ( .A(n36), .Z(n41) );
  BUF_X1 U10 ( .A(n37), .Z(n46) );
  BUF_X1 U11 ( .A(n38), .Z(n48) );
  BUF_X1 U12 ( .A(n36), .Z(n42) );
  BUF_X1 U13 ( .A(n36), .Z(n43) );
  BUF_X1 U14 ( .A(n37), .Z(n45) );
  BUF_X1 U15 ( .A(n38), .Z(n47) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n36) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n37) );
  OAI22_X1 U19 ( .A1(n69), .A2(n40), .B1(n41), .B2(n56), .ZN(n7) );
  INV_X1 U20 ( .A(D[28]), .ZN(n56) );
  OAI22_X1 U21 ( .A1(n70), .A2(n39), .B1(n41), .B2(n57), .ZN(n8) );
  INV_X1 U22 ( .A(D[27]), .ZN(n57) );
  OAI22_X1 U23 ( .A1(n68), .A2(n40), .B1(n41), .B2(n55), .ZN(n6) );
  INV_X1 U24 ( .A(D[29]), .ZN(n55) );
  OAI22_X1 U25 ( .A1(n96), .A2(n39), .B1(n42), .B2(n115), .ZN(n34) );
  INV_X1 U26 ( .A(D[1]), .ZN(n115) );
  OAI22_X1 U27 ( .A1(n97), .A2(n39), .B1(n42), .B2(n116), .ZN(n35) );
  INV_X1 U28 ( .A(D[0]), .ZN(n116) );
  OAI22_X1 U29 ( .A1(n71), .A2(n40), .B1(n41), .B2(n58), .ZN(n9) );
  INV_X1 U30 ( .A(D[26]), .ZN(n58) );
  OAI22_X1 U31 ( .A1(n67), .A2(n39), .B1(n42), .B2(n54), .ZN(n5) );
  INV_X1 U32 ( .A(D[30]), .ZN(n54) );
  OAI22_X1 U33 ( .A1(n66), .A2(n40), .B1(n42), .B2(n53), .ZN(n4) );
  INV_X1 U34 ( .A(D[31]), .ZN(n53) );
  OAI22_X1 U35 ( .A1(n85), .A2(n40), .B1(n45), .B2(n104), .ZN(n23) );
  INV_X1 U36 ( .A(D[12]), .ZN(n104) );
  OAI22_X1 U37 ( .A1(n84), .A2(n40), .B1(n45), .B2(n103), .ZN(n22) );
  INV_X1 U38 ( .A(D[13]), .ZN(n103) );
  OAI22_X1 U39 ( .A1(n90), .A2(n40), .B1(n44), .B2(n109), .ZN(n28) );
  INV_X1 U40 ( .A(D[7]), .ZN(n109) );
  OAI22_X1 U41 ( .A1(n87), .A2(n40), .B1(n45), .B2(n106), .ZN(n25) );
  INV_X1 U42 ( .A(D[10]), .ZN(n106) );
  OAI22_X1 U43 ( .A1(n77), .A2(n39), .B1(n47), .B2(n64), .ZN(n15) );
  INV_X1 U44 ( .A(D[20]), .ZN(n64) );
  OAI22_X1 U45 ( .A1(n91), .A2(n40), .B1(n44), .B2(n110), .ZN(n29) );
  INV_X1 U46 ( .A(D[6]), .ZN(n110) );
  OAI22_X1 U47 ( .A1(n93), .A2(n40), .B1(n43), .B2(n112), .ZN(n31) );
  INV_X1 U48 ( .A(D[4]), .ZN(n112) );
  OAI22_X1 U49 ( .A1(n80), .A2(n39), .B1(n46), .B2(n99), .ZN(n18) );
  INV_X1 U50 ( .A(D[17]), .ZN(n99) );
  OAI22_X1 U51 ( .A1(n88), .A2(n40), .B1(n44), .B2(n107), .ZN(n26) );
  INV_X1 U52 ( .A(D[9]), .ZN(n107) );
  OAI22_X1 U53 ( .A1(n83), .A2(n39), .B1(n46), .B2(n102), .ZN(n21) );
  INV_X1 U54 ( .A(D[14]), .ZN(n102) );
  OAI22_X1 U55 ( .A1(n89), .A2(n40), .B1(n44), .B2(n108), .ZN(n27) );
  INV_X1 U56 ( .A(D[8]), .ZN(n108) );
  OAI22_X1 U57 ( .A1(n72), .A2(n39), .B1(n48), .B2(n59), .ZN(n10) );
  INV_X1 U58 ( .A(D[25]), .ZN(n59) );
  OAI22_X1 U59 ( .A1(n92), .A2(n40), .B1(n43), .B2(n111), .ZN(n30) );
  INV_X1 U60 ( .A(D[5]), .ZN(n111) );
  OAI22_X1 U61 ( .A1(n82), .A2(n39), .B1(n46), .B2(n101), .ZN(n20) );
  INV_X1 U62 ( .A(D[15]), .ZN(n101) );
  OAI22_X1 U63 ( .A1(n81), .A2(n39), .B1(n46), .B2(n100), .ZN(n19) );
  INV_X1 U64 ( .A(D[16]), .ZN(n100) );
  OAI22_X1 U65 ( .A1(n76), .A2(n39), .B1(n47), .B2(n63), .ZN(n14) );
  INV_X1 U66 ( .A(D[21]), .ZN(n63) );
  OAI22_X1 U67 ( .A1(n75), .A2(n39), .B1(n48), .B2(n62), .ZN(n13) );
  INV_X1 U68 ( .A(D[22]), .ZN(n62) );
  OAI22_X1 U69 ( .A1(n73), .A2(n39), .B1(n48), .B2(n60), .ZN(n11) );
  INV_X1 U70 ( .A(D[24]), .ZN(n60) );
  OAI22_X1 U71 ( .A1(n74), .A2(n39), .B1(n48), .B2(n61), .ZN(n12) );
  INV_X1 U72 ( .A(D[23]), .ZN(n61) );
  OAI22_X1 U73 ( .A1(n95), .A2(n40), .B1(n43), .B2(n114), .ZN(n33) );
  INV_X1 U74 ( .A(D[2]), .ZN(n114) );
  OAI22_X1 U75 ( .A1(n94), .A2(n40), .B1(n43), .B2(n113), .ZN(n32) );
  INV_X1 U76 ( .A(D[3]), .ZN(n113) );
  OAI22_X1 U77 ( .A1(n86), .A2(n40), .B1(n45), .B2(n105), .ZN(n24) );
  INV_X1 U78 ( .A(D[11]), .ZN(n105) );
  OAI22_X1 U79 ( .A1(n79), .A2(n39), .B1(n47), .B2(n98), .ZN(n17) );
  INV_X1 U80 ( .A(D[18]), .ZN(n98) );
  OAI22_X1 U81 ( .A1(n78), .A2(n39), .B1(n47), .B2(n65), .ZN(n16) );
  INV_X1 U82 ( .A(D[19]), .ZN(n65) );
endmodule


module REG_GEN_NBIT32_11 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n52), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n52), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n52), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n52), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n52), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n51), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n51), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n51), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n51), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n51), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n51), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n52), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n52), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n50), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n50), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n50), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n50), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n50), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n50), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n50), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n50), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n50), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n50), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n50), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n50), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n51), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n52), .Q(Q[0]), .QN(n97) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n45) );
  BUF_X1 U10 ( .A(n37), .Z(n46) );
  BUF_X1 U11 ( .A(n36), .Z(n42) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n37), .Z(n44) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n71), .A2(n40), .B1(n41), .B2(n58), .ZN(n9) );
  INV_X1 U20 ( .A(D[26]), .ZN(n58) );
  OAI22_X1 U21 ( .A1(n70), .A2(n39), .B1(n41), .B2(n57), .ZN(n8) );
  INV_X1 U22 ( .A(D[27]), .ZN(n57) );
  OAI22_X1 U23 ( .A1(n68), .A2(n40), .B1(n41), .B2(n55), .ZN(n6) );
  INV_X1 U24 ( .A(D[29]), .ZN(n55) );
  OAI22_X1 U25 ( .A1(n67), .A2(n39), .B1(n42), .B2(n54), .ZN(n5) );
  INV_X1 U26 ( .A(D[30]), .ZN(n54) );
  OAI22_X1 U27 ( .A1(n66), .A2(n40), .B1(n42), .B2(n53), .ZN(n4) );
  INV_X1 U28 ( .A(D[31]), .ZN(n53) );
  OAI22_X1 U29 ( .A1(n97), .A2(n39), .B1(n42), .B2(n116), .ZN(n35) );
  INV_X1 U30 ( .A(D[0]), .ZN(n116) );
  OAI22_X1 U31 ( .A1(n96), .A2(n40), .B1(n42), .B2(n115), .ZN(n34) );
  INV_X1 U32 ( .A(D[1]), .ZN(n115) );
  INV_X1 U33 ( .A(D[6]), .ZN(n110) );
  INV_X1 U34 ( .A(D[8]), .ZN(n108) );
  INV_X1 U35 ( .A(D[21]), .ZN(n63) );
  INV_X1 U36 ( .A(D[22]), .ZN(n62) );
  INV_X1 U37 ( .A(D[28]), .ZN(n56) );
  OAI22_X1 U38 ( .A1(n95), .A2(n40), .B1(n43), .B2(n114), .ZN(n33) );
  INV_X1 U39 ( .A(D[2]), .ZN(n114) );
  OAI22_X1 U40 ( .A1(n94), .A2(n40), .B1(n43), .B2(n113), .ZN(n32) );
  INV_X1 U41 ( .A(D[3]), .ZN(n113) );
  OAI22_X1 U42 ( .A1(n93), .A2(n40), .B1(n43), .B2(n112), .ZN(n31) );
  INV_X1 U43 ( .A(D[4]), .ZN(n112) );
  OAI22_X1 U44 ( .A1(n92), .A2(n40), .B1(n43), .B2(n111), .ZN(n30) );
  INV_X1 U45 ( .A(D[5]), .ZN(n111) );
  OAI22_X1 U46 ( .A1(n90), .A2(n40), .B1(n44), .B2(n109), .ZN(n28) );
  INV_X1 U47 ( .A(D[7]), .ZN(n109) );
  OAI22_X1 U48 ( .A1(n88), .A2(n40), .B1(n44), .B2(n107), .ZN(n26) );
  INV_X1 U49 ( .A(D[9]), .ZN(n107) );
  OAI22_X1 U50 ( .A1(n87), .A2(n40), .B1(n45), .B2(n106), .ZN(n25) );
  INV_X1 U51 ( .A(D[10]), .ZN(n106) );
  OAI22_X1 U52 ( .A1(n86), .A2(n40), .B1(n45), .B2(n105), .ZN(n24) );
  INV_X1 U53 ( .A(D[11]), .ZN(n105) );
  OAI22_X1 U54 ( .A1(n85), .A2(n40), .B1(n45), .B2(n104), .ZN(n23) );
  INV_X1 U55 ( .A(D[12]), .ZN(n104) );
  OAI22_X1 U56 ( .A1(n84), .A2(n40), .B1(n45), .B2(n103), .ZN(n22) );
  INV_X1 U57 ( .A(D[13]), .ZN(n103) );
  OAI22_X1 U58 ( .A1(n83), .A2(n39), .B1(n46), .B2(n102), .ZN(n21) );
  INV_X1 U59 ( .A(D[14]), .ZN(n102) );
  OAI22_X1 U60 ( .A1(n82), .A2(n39), .B1(n46), .B2(n101), .ZN(n20) );
  INV_X1 U61 ( .A(D[15]), .ZN(n101) );
  OAI22_X1 U62 ( .A1(n81), .A2(n39), .B1(n46), .B2(n100), .ZN(n19) );
  INV_X1 U63 ( .A(D[16]), .ZN(n100) );
  OAI22_X1 U64 ( .A1(n80), .A2(n39), .B1(n46), .B2(n99), .ZN(n18) );
  INV_X1 U65 ( .A(D[17]), .ZN(n99) );
  OAI22_X1 U66 ( .A1(n79), .A2(n39), .B1(n47), .B2(n98), .ZN(n17) );
  INV_X1 U67 ( .A(D[18]), .ZN(n98) );
  OAI22_X1 U68 ( .A1(n78), .A2(n39), .B1(n47), .B2(n65), .ZN(n16) );
  INV_X1 U69 ( .A(D[19]), .ZN(n65) );
  OAI22_X1 U70 ( .A1(n77), .A2(n39), .B1(n47), .B2(n64), .ZN(n15) );
  INV_X1 U71 ( .A(D[20]), .ZN(n64) );
  OAI22_X1 U72 ( .A1(n74), .A2(n39), .B1(n48), .B2(n61), .ZN(n12) );
  INV_X1 U73 ( .A(D[23]), .ZN(n61) );
  OAI22_X1 U74 ( .A1(n73), .A2(n39), .B1(n48), .B2(n60), .ZN(n11) );
  INV_X1 U75 ( .A(D[24]), .ZN(n60) );
  OAI22_X1 U76 ( .A1(n72), .A2(n39), .B1(n48), .B2(n59), .ZN(n10) );
  INV_X1 U77 ( .A(D[25]), .ZN(n59) );
  OAI22_X1 U78 ( .A1(n69), .A2(n39), .B1(n41), .B2(n56), .ZN(n7) );
  OAI22_X1 U79 ( .A1(n91), .A2(n40), .B1(n44), .B2(n110), .ZN(n29) );
  OAI22_X1 U80 ( .A1(n76), .A2(n39), .B1(n47), .B2(n63), .ZN(n14) );
  OAI22_X1 U81 ( .A1(n75), .A2(n39), .B1(n48), .B2(n62), .ZN(n13) );
  OAI22_X1 U82 ( .A1(n89), .A2(n40), .B1(n44), .B2(n108), .ZN(n27) );
endmodule


module REG_GEN_NBIT32_10 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n50), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n50), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n50), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n50), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n50), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n50), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n50), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n50), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n50), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n50), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n50), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n50), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n51), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n51), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n51), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n51), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n51), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n51), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n51), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n52), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n52), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n52), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n52), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n52), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n52), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n52), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n52), .Q(Q[0]), .QN(n97) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n44) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n97), .A2(n40), .B1(n42), .B2(n116), .ZN(n35) );
  INV_X1 U20 ( .A(D[0]), .ZN(n116) );
  OAI22_X1 U21 ( .A1(n96), .A2(n39), .B1(n42), .B2(n115), .ZN(n34) );
  INV_X1 U22 ( .A(D[1]), .ZN(n115) );
  OAI22_X1 U23 ( .A1(n71), .A2(n40), .B1(n41), .B2(n58), .ZN(n9) );
  INV_X1 U24 ( .A(D[26]), .ZN(n58) );
  OAI22_X1 U25 ( .A1(n70), .A2(n39), .B1(n41), .B2(n57), .ZN(n8) );
  INV_X1 U26 ( .A(D[27]), .ZN(n57) );
  OAI22_X1 U27 ( .A1(n69), .A2(n40), .B1(n41), .B2(n56), .ZN(n7) );
  INV_X1 U28 ( .A(D[28]), .ZN(n56) );
  OAI22_X1 U29 ( .A1(n68), .A2(n39), .B1(n41), .B2(n55), .ZN(n6) );
  INV_X1 U30 ( .A(D[29]), .ZN(n55) );
  OAI22_X1 U31 ( .A1(n67), .A2(n40), .B1(n42), .B2(n54), .ZN(n5) );
  INV_X1 U32 ( .A(D[30]), .ZN(n54) );
  OAI22_X1 U33 ( .A1(n66), .A2(n39), .B1(n42), .B2(n53), .ZN(n4) );
  INV_X1 U34 ( .A(D[31]), .ZN(n53) );
  OAI22_X1 U35 ( .A1(n95), .A2(n40), .B1(n43), .B2(n114), .ZN(n33) );
  INV_X1 U36 ( .A(D[2]), .ZN(n114) );
  OAI22_X1 U37 ( .A1(n94), .A2(n40), .B1(n43), .B2(n113), .ZN(n32) );
  INV_X1 U38 ( .A(D[3]), .ZN(n113) );
  OAI22_X1 U39 ( .A1(n93), .A2(n40), .B1(n43), .B2(n112), .ZN(n31) );
  INV_X1 U40 ( .A(D[4]), .ZN(n112) );
  OAI22_X1 U41 ( .A1(n92), .A2(n40), .B1(n43), .B2(n111), .ZN(n30) );
  INV_X1 U42 ( .A(D[5]), .ZN(n111) );
  OAI22_X1 U43 ( .A1(n91), .A2(n40), .B1(n44), .B2(n110), .ZN(n29) );
  INV_X1 U44 ( .A(D[6]), .ZN(n110) );
  OAI22_X1 U45 ( .A1(n90), .A2(n40), .B1(n44), .B2(n109), .ZN(n28) );
  INV_X1 U46 ( .A(D[7]), .ZN(n109) );
  OAI22_X1 U47 ( .A1(n89), .A2(n40), .B1(n44), .B2(n108), .ZN(n27) );
  INV_X1 U48 ( .A(D[8]), .ZN(n108) );
  OAI22_X1 U49 ( .A1(n88), .A2(n40), .B1(n44), .B2(n107), .ZN(n26) );
  INV_X1 U50 ( .A(D[9]), .ZN(n107) );
  OAI22_X1 U51 ( .A1(n87), .A2(n40), .B1(n45), .B2(n106), .ZN(n25) );
  INV_X1 U52 ( .A(D[10]), .ZN(n106) );
  OAI22_X1 U53 ( .A1(n86), .A2(n40), .B1(n45), .B2(n105), .ZN(n24) );
  INV_X1 U54 ( .A(D[11]), .ZN(n105) );
  OAI22_X1 U55 ( .A1(n85), .A2(n40), .B1(n45), .B2(n104), .ZN(n23) );
  INV_X1 U56 ( .A(D[12]), .ZN(n104) );
  OAI22_X1 U57 ( .A1(n84), .A2(n40), .B1(n45), .B2(n103), .ZN(n22) );
  INV_X1 U58 ( .A(D[13]), .ZN(n103) );
  OAI22_X1 U59 ( .A1(n83), .A2(n39), .B1(n46), .B2(n102), .ZN(n21) );
  INV_X1 U60 ( .A(D[14]), .ZN(n102) );
  OAI22_X1 U61 ( .A1(n82), .A2(n39), .B1(n46), .B2(n101), .ZN(n20) );
  INV_X1 U62 ( .A(D[15]), .ZN(n101) );
  OAI22_X1 U63 ( .A1(n81), .A2(n39), .B1(n46), .B2(n100), .ZN(n19) );
  INV_X1 U64 ( .A(D[16]), .ZN(n100) );
  OAI22_X1 U65 ( .A1(n80), .A2(n39), .B1(n46), .B2(n99), .ZN(n18) );
  INV_X1 U66 ( .A(D[17]), .ZN(n99) );
  OAI22_X1 U67 ( .A1(n79), .A2(n39), .B1(n47), .B2(n98), .ZN(n17) );
  INV_X1 U68 ( .A(D[18]), .ZN(n98) );
  OAI22_X1 U69 ( .A1(n78), .A2(n39), .B1(n47), .B2(n65), .ZN(n16) );
  INV_X1 U70 ( .A(D[19]), .ZN(n65) );
  OAI22_X1 U71 ( .A1(n77), .A2(n39), .B1(n47), .B2(n64), .ZN(n15) );
  INV_X1 U72 ( .A(D[20]), .ZN(n64) );
  OAI22_X1 U73 ( .A1(n76), .A2(n39), .B1(n47), .B2(n63), .ZN(n14) );
  INV_X1 U74 ( .A(D[21]), .ZN(n63) );
  OAI22_X1 U75 ( .A1(n75), .A2(n39), .B1(n48), .B2(n62), .ZN(n13) );
  INV_X1 U76 ( .A(D[22]), .ZN(n62) );
  OAI22_X1 U77 ( .A1(n74), .A2(n39), .B1(n48), .B2(n61), .ZN(n12) );
  INV_X1 U78 ( .A(D[23]), .ZN(n61) );
  OAI22_X1 U79 ( .A1(n73), .A2(n39), .B1(n48), .B2(n60), .ZN(n11) );
  INV_X1 U80 ( .A(D[24]), .ZN(n60) );
  OAI22_X1 U81 ( .A1(n72), .A2(n39), .B1(n48), .B2(n59), .ZN(n10) );
  INV_X1 U82 ( .A(D[25]), .ZN(n59) );
endmodule


module decodeUnit_nbit32 ( Clk, Rst, en_reg, RD1, RD2, IRAM_instr, PC_Next, WR, 
        ADD_RW, DATA_RW, RW_R_out, RW_I_out, Jump_address, I_immediate_ext_out, 
        RD_data_1_out, RD_data_2_out, PC_Next_out, Opcode, Func );
  input [31:0] IRAM_instr;
  input [31:0] PC_Next;
  input [4:0] ADD_RW;
  input [31:0] DATA_RW;
  output [31:0] RW_R_out;
  output [31:0] RW_I_out;
  output [31:0] Jump_address;
  output [31:0] I_immediate_ext_out;
  output [31:0] RD_data_1_out;
  output [31:0] RD_data_2_out;
  output [31:0] PC_Next_out;
  output [5:0] Opcode;
  output [10:0] Func;
  input Clk, Rst, en_reg, RD1, RD2, WR;
  wire   \IRAM_instr[31] , \IRAM_instr[30] , \IRAM_instr[29] ,
         \IRAM_instr[28] , \IRAM_instr[27] , \IRAM_instr[26] ,
         \IRAM_instr[10] , \IRAM_instr[9] , \IRAM_instr[8] , \IRAM_instr[7] ,
         \IRAM_instr[6] , \IRAM_instr[5] , \IRAM_instr[4] , \IRAM_instr[3] ,
         \IRAM_instr[2] , \IRAM_instr[1] , \IRAM_instr[0] , n1;
  wire   [31:0] Jump_addr;
  wire   [31:0] RD_data_1;
  wire   [31:0] RD_data_2;
  wire   [31:0] I_immediate_ext;
  assign Opcode[5] = \IRAM_instr[31] ;
  assign \IRAM_instr[31]  = IRAM_instr[31];
  assign Opcode[4] = \IRAM_instr[30] ;
  assign \IRAM_instr[30]  = IRAM_instr[30];
  assign Opcode[3] = \IRAM_instr[29] ;
  assign \IRAM_instr[29]  = IRAM_instr[29];
  assign Opcode[2] = \IRAM_instr[28] ;
  assign \IRAM_instr[28]  = IRAM_instr[28];
  assign Opcode[1] = \IRAM_instr[27] ;
  assign \IRAM_instr[27]  = IRAM_instr[27];
  assign Opcode[0] = \IRAM_instr[26] ;
  assign \IRAM_instr[26]  = IRAM_instr[26];
  assign Func[10] = \IRAM_instr[10] ;
  assign \IRAM_instr[10]  = IRAM_instr[10];
  assign Func[9] = \IRAM_instr[9] ;
  assign \IRAM_instr[9]  = IRAM_instr[9];
  assign Func[8] = \IRAM_instr[8] ;
  assign \IRAM_instr[8]  = IRAM_instr[8];
  assign Func[7] = \IRAM_instr[7] ;
  assign \IRAM_instr[7]  = IRAM_instr[7];
  assign Func[6] = \IRAM_instr[6] ;
  assign \IRAM_instr[6]  = IRAM_instr[6];
  assign Func[5] = \IRAM_instr[5] ;
  assign \IRAM_instr[5]  = IRAM_instr[5];
  assign Func[4] = \IRAM_instr[4] ;
  assign \IRAM_instr[4]  = IRAM_instr[4];
  assign Func[3] = \IRAM_instr[3] ;
  assign \IRAM_instr[3]  = IRAM_instr[3];
  assign Func[2] = \IRAM_instr[2] ;
  assign \IRAM_instr[2]  = IRAM_instr[2];
  assign Func[1] = \IRAM_instr[1] ;
  assign \IRAM_instr[1]  = IRAM_instr[1];
  assign Func[0] = \IRAM_instr[0] ;
  assign \IRAM_instr[0]  = IRAM_instr[0];

  sign_extension_sign_init26_sign_ext32 SIGN_EXT_immediate_J ( .data_in({
        IRAM_instr[25:11], \IRAM_instr[10] , \IRAM_instr[9] , \IRAM_instr[8] , 
        \IRAM_instr[7] , \IRAM_instr[6] , \IRAM_instr[5] , \IRAM_instr[4] , 
        \IRAM_instr[3] , \IRAM_instr[2] , \IRAM_instr[1] , \IRAM_instr[0] }), 
        .data_out(Jump_addr) );
  register_file_nbit_reg32_n_reg32_nbit_addr5 REGISTERS ( .reset(Rst), 
        .enable(1'b0), .rd1(RD1), .rd2(RD2), .wr(WR), .add_wr(ADD_RW), 
        .add_rd1(IRAM_instr[25:21]), .add_rd2(IRAM_instr[20:16]), .datain(
        DATA_RW), .out1(RD_data_1), .out2(RD_data_2) );
  sign_extension_sign_init16_sign_ext32 SIGN_EXT_immediate_I ( .data_in({
        IRAM_instr[15:11], \IRAM_instr[10] , \IRAM_instr[9] , \IRAM_instr[8] , 
        \IRAM_instr[7] , \IRAM_instr[6] , \IRAM_instr[5] , \IRAM_instr[4] , 
        \IRAM_instr[3] , \IRAM_instr[2] , \IRAM_instr[1] , \IRAM_instr[0] }), 
        .data_out(I_immediate_ext) );
  REG_GEN_NBIT32_16 ID_reg_RW_R ( .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, IRAM_instr[15:11]}), 
        .CK(Clk), .Enable_n(n1), .RESET_n(Rst), .Q(RW_R_out) );
  REG_GEN_NBIT32_15 ID_reg_RW_I ( .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, IRAM_instr[20:16]}), 
        .CK(Clk), .Enable_n(n1), .RESET_n(Rst), .Q(RW_I_out) );
  REG_GEN_NBIT32_14 ID_reg_I_imm ( .D(I_immediate_ext), .CK(Clk), .Enable_n(n1), .RESET_n(Rst), .Q(I_immediate_ext_out) );
  REG_GEN_NBIT32_13 ID_reg_J_imm ( .D(Jump_addr), .CK(Clk), .Enable_n(n1), 
        .RESET_n(Rst), .Q(Jump_address) );
  REG_GEN_NBIT32_12 ID_reg_RD_data_1 ( .D(RD_data_1), .CK(Clk), .Enable_n(n1), 
        .RESET_n(Rst), .Q(RD_data_1_out) );
  REG_GEN_NBIT32_11 ID_reg_RD_data_2 ( .D(RD_data_2), .CK(Clk), .Enable_n(n1), 
        .RESET_n(Rst), .Q(RD_data_2_out) );
  REG_GEN_NBIT32_10 ID_reg_PC_next ( .D(PC_Next), .CK(Clk), .Enable_n(n1), 
        .RESET_n(Rst), .Q(PC_Next_out) );
  BUF_X1 U2 ( .A(en_reg), .Z(n1) );
endmodule


module MUX21_GENERIC_NBIT32_8 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n33, n66, n67, n100;

  INV_X1 U1 ( .A(n39), .ZN(Y[4]) );
  INV_X1 U2 ( .A(n58), .ZN(Y[16]) );
  INV_X1 U3 ( .A(n57), .ZN(Y[17]) );
  INV_X1 U4 ( .A(n56), .ZN(Y[18]) );
  INV_X1 U5 ( .A(n48), .ZN(Y[25]) );
  INV_X1 U6 ( .A(n46), .ZN(Y[27]) );
  INV_X1 U7 ( .A(n42), .ZN(Y[30]) );
  INV_X1 U8 ( .A(n64), .ZN(Y[10]) );
  INV_X1 U9 ( .A(n62), .ZN(Y[12]) );
  INV_X1 U10 ( .A(n63), .ZN(Y[11]) );
  INV_X1 U11 ( .A(n38), .ZN(Y[5]) );
  INV_X1 U12 ( .A(n40), .ZN(Y[3]) );
  INV_X1 U13 ( .A(n50), .ZN(Y[23]) );
  BUF_X1 U14 ( .A(n100), .Z(n33) );
  BUF_X1 U15 ( .A(n100), .Z(n66) );
  BUF_X1 U16 ( .A(n100), .Z(n67) );
  AOI22_X1 U17 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(SEL), .ZN(n40) );
  AOI22_X1 U18 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(SEL), .ZN(n39) );
  AOI22_X1 U19 ( .A1(A[11]), .A2(n33), .B1(B[11]), .B2(SEL), .ZN(n63) );
  AOI22_X1 U20 ( .A1(A[12]), .A2(n33), .B1(B[12]), .B2(SEL), .ZN(n62) );
  AOI22_X1 U21 ( .A1(A[10]), .A2(n33), .B1(B[10]), .B2(SEL), .ZN(n64) );
  AOI22_X1 U22 ( .A1(A[17]), .A2(n33), .B1(B[17]), .B2(SEL), .ZN(n57) );
  AOI22_X1 U23 ( .A1(A[16]), .A2(n33), .B1(B[16]), .B2(SEL), .ZN(n58) );
  AOI22_X1 U24 ( .A1(A[18]), .A2(n33), .B1(B[18]), .B2(SEL), .ZN(n56) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(SEL), .ZN(n38) );
  AOI22_X1 U26 ( .A1(A[30]), .A2(n66), .B1(B[30]), .B2(SEL), .ZN(n42) );
  AOI22_X1 U27 ( .A1(A[27]), .A2(n66), .B1(B[27]), .B2(SEL), .ZN(n46) );
  AOI22_X1 U28 ( .A1(A[23]), .A2(n66), .B1(B[23]), .B2(SEL), .ZN(n50) );
  AOI22_X1 U29 ( .A1(A[25]), .A2(n66), .B1(B[25]), .B2(SEL), .ZN(n48) );
  INV_X1 U30 ( .A(n59), .ZN(Y[15]) );
  AOI22_X1 U31 ( .A1(A[15]), .A2(n33), .B1(B[15]), .B2(SEL), .ZN(n59) );
  INV_X1 U32 ( .A(n53), .ZN(Y[20]) );
  AOI22_X1 U33 ( .A1(A[20]), .A2(n66), .B1(B[20]), .B2(SEL), .ZN(n53) );
  INV_X1 U34 ( .A(n49), .ZN(Y[24]) );
  AOI22_X1 U35 ( .A1(A[24]), .A2(n66), .B1(B[24]), .B2(SEL), .ZN(n49) );
  INV_X1 U36 ( .A(n41), .ZN(Y[31]) );
  AOI22_X1 U37 ( .A1(A[31]), .A2(n67), .B1(B[31]), .B2(SEL), .ZN(n41) );
  INV_X1 U38 ( .A(n60), .ZN(Y[14]) );
  AOI22_X1 U39 ( .A1(A[14]), .A2(n33), .B1(B[14]), .B2(SEL), .ZN(n60) );
  INV_X1 U40 ( .A(n61), .ZN(Y[13]) );
  AOI22_X1 U41 ( .A1(A[13]), .A2(n33), .B1(B[13]), .B2(SEL), .ZN(n61) );
  INV_X1 U42 ( .A(n36), .ZN(Y[7]) );
  AOI22_X1 U43 ( .A1(A[7]), .A2(n67), .B1(B[7]), .B2(SEL), .ZN(n36) );
  AOI22_X1 U44 ( .A1(A[9]), .A2(n67), .B1(SEL), .B2(B[9]), .ZN(n34) );
  AOI22_X1 U45 ( .A1(A[2]), .A2(n66), .B1(B[2]), .B2(SEL), .ZN(n43) );
  AOI22_X1 U46 ( .A1(A[1]), .A2(n33), .B1(B[1]), .B2(SEL), .ZN(n54) );
  AOI22_X1 U47 ( .A1(A[0]), .A2(n33), .B1(B[0]), .B2(SEL), .ZN(n65) );
  INV_X1 U48 ( .A(SEL), .ZN(n100) );
  INV_X1 U49 ( .A(n54), .ZN(Y[1]) );
  INV_X1 U50 ( .A(n43), .ZN(Y[2]) );
  INV_X1 U51 ( .A(n65), .ZN(Y[0]) );
  INV_X1 U52 ( .A(n55), .ZN(Y[19]) );
  AOI22_X1 U53 ( .A1(A[26]), .A2(n66), .B1(B[26]), .B2(SEL), .ZN(n47) );
  INV_X1 U54 ( .A(n47), .ZN(Y[26]) );
  AOI22_X1 U55 ( .A1(A[19]), .A2(n33), .B1(B[19]), .B2(SEL), .ZN(n55) );
  INV_X1 U56 ( .A(n37), .ZN(Y[6]) );
  AOI22_X1 U57 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(SEL), .ZN(n37) );
  INV_X1 U58 ( .A(n34), .ZN(Y[9]) );
  INV_X1 U59 ( .A(n51), .ZN(Y[22]) );
  AOI22_X1 U60 ( .A1(A[22]), .A2(n66), .B1(B[22]), .B2(SEL), .ZN(n51) );
  INV_X1 U61 ( .A(n44), .ZN(Y[29]) );
  AOI22_X1 U62 ( .A1(A[29]), .A2(n66), .B1(B[29]), .B2(SEL), .ZN(n44) );
  AOI22_X1 U63 ( .A1(A[8]), .A2(n67), .B1(B[8]), .B2(SEL), .ZN(n35) );
  INV_X1 U64 ( .A(n35), .ZN(Y[8]) );
  INV_X1 U65 ( .A(n45), .ZN(Y[28]) );
  AOI22_X1 U66 ( .A1(A[28]), .A2(n66), .B1(B[28]), .B2(SEL), .ZN(n45) );
  AOI22_X1 U67 ( .A1(A[21]), .A2(n66), .B1(B[21]), .B2(SEL), .ZN(n52) );
  INV_X1 U68 ( .A(n52), .ZN(Y[21]) );
endmodule


module MUX21_GENERIC_NBIT32_7 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n33, n66, n67, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132;

  BUF_X1 U1 ( .A(n100), .Z(n33) );
  BUF_X1 U2 ( .A(n100), .Z(n66) );
  BUF_X1 U3 ( .A(n100), .Z(n67) );
  INV_X1 U4 ( .A(n101), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n33), .B1(B[0]), .B2(SEL), .ZN(n101) );
  INV_X1 U6 ( .A(n112), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n33), .B1(B[1]), .B2(SEL), .ZN(n112) );
  INV_X1 U8 ( .A(n119), .ZN(Y[26]) );
  AOI22_X1 U9 ( .A1(A[26]), .A2(n66), .B1(B[26]), .B2(SEL), .ZN(n119) );
  INV_X1 U10 ( .A(n120), .ZN(Y[27]) );
  AOI22_X1 U11 ( .A1(A[27]), .A2(n66), .B1(B[27]), .B2(SEL), .ZN(n120) );
  INV_X1 U12 ( .A(n121), .ZN(Y[28]) );
  AOI22_X1 U13 ( .A1(A[28]), .A2(n66), .B1(B[28]), .B2(SEL), .ZN(n121) );
  INV_X1 U14 ( .A(n122), .ZN(Y[29]) );
  AOI22_X1 U15 ( .A1(A[29]), .A2(n66), .B1(B[29]), .B2(SEL), .ZN(n122) );
  INV_X1 U16 ( .A(n124), .ZN(Y[30]) );
  AOI22_X1 U17 ( .A1(A[30]), .A2(n66), .B1(B[30]), .B2(SEL), .ZN(n124) );
  INV_X1 U18 ( .A(n125), .ZN(Y[31]) );
  AOI22_X1 U19 ( .A1(A[31]), .A2(n67), .B1(B[31]), .B2(SEL), .ZN(n125) );
  INV_X1 U20 ( .A(n104), .ZN(Y[12]) );
  AOI22_X1 U21 ( .A1(A[12]), .A2(n33), .B1(B[12]), .B2(SEL), .ZN(n104) );
  INV_X1 U22 ( .A(n105), .ZN(Y[13]) );
  AOI22_X1 U23 ( .A1(A[13]), .A2(n33), .B1(B[13]), .B2(SEL), .ZN(n105) );
  INV_X1 U24 ( .A(n106), .ZN(Y[14]) );
  AOI22_X1 U25 ( .A1(A[14]), .A2(n33), .B1(B[14]), .B2(SEL), .ZN(n106) );
  INV_X1 U26 ( .A(n107), .ZN(Y[15]) );
  AOI22_X1 U27 ( .A1(A[15]), .A2(n33), .B1(B[15]), .B2(SEL), .ZN(n107) );
  INV_X1 U28 ( .A(n108), .ZN(Y[16]) );
  AOI22_X1 U29 ( .A1(A[16]), .A2(n33), .B1(B[16]), .B2(SEL), .ZN(n108) );
  INV_X1 U30 ( .A(n109), .ZN(Y[17]) );
  AOI22_X1 U31 ( .A1(A[17]), .A2(n33), .B1(B[17]), .B2(SEL), .ZN(n109) );
  INV_X1 U32 ( .A(n110), .ZN(Y[18]) );
  AOI22_X1 U33 ( .A1(A[18]), .A2(n33), .B1(B[18]), .B2(SEL), .ZN(n110) );
  INV_X1 U34 ( .A(n111), .ZN(Y[19]) );
  AOI22_X1 U35 ( .A1(A[19]), .A2(n33), .B1(B[19]), .B2(SEL), .ZN(n111) );
  INV_X1 U36 ( .A(n113), .ZN(Y[20]) );
  AOI22_X1 U37 ( .A1(A[20]), .A2(n66), .B1(B[20]), .B2(SEL), .ZN(n113) );
  INV_X1 U38 ( .A(n114), .ZN(Y[21]) );
  AOI22_X1 U39 ( .A1(A[21]), .A2(n66), .B1(B[21]), .B2(SEL), .ZN(n114) );
  INV_X1 U40 ( .A(n115), .ZN(Y[22]) );
  AOI22_X1 U41 ( .A1(A[22]), .A2(n66), .B1(B[22]), .B2(SEL), .ZN(n115) );
  INV_X1 U42 ( .A(n116), .ZN(Y[23]) );
  AOI22_X1 U43 ( .A1(A[23]), .A2(n66), .B1(B[23]), .B2(SEL), .ZN(n116) );
  INV_X1 U44 ( .A(n117), .ZN(Y[24]) );
  AOI22_X1 U45 ( .A1(A[24]), .A2(n66), .B1(B[24]), .B2(SEL), .ZN(n117) );
  INV_X1 U46 ( .A(n118), .ZN(Y[25]) );
  AOI22_X1 U47 ( .A1(A[25]), .A2(n66), .B1(B[25]), .B2(SEL), .ZN(n118) );
  INV_X1 U48 ( .A(n123), .ZN(Y[2]) );
  AOI22_X1 U49 ( .A1(A[2]), .A2(n66), .B1(B[2]), .B2(SEL), .ZN(n123) );
  INV_X1 U50 ( .A(n126), .ZN(Y[3]) );
  AOI22_X1 U51 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(SEL), .ZN(n126) );
  INV_X1 U52 ( .A(n127), .ZN(Y[4]) );
  AOI22_X1 U53 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(SEL), .ZN(n127) );
  INV_X1 U54 ( .A(n128), .ZN(Y[5]) );
  AOI22_X1 U55 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(SEL), .ZN(n128) );
  INV_X1 U56 ( .A(n129), .ZN(Y[6]) );
  AOI22_X1 U57 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(SEL), .ZN(n129) );
  INV_X1 U58 ( .A(n130), .ZN(Y[7]) );
  AOI22_X1 U59 ( .A1(A[7]), .A2(n67), .B1(B[7]), .B2(SEL), .ZN(n130) );
  INV_X1 U60 ( .A(n131), .ZN(Y[8]) );
  AOI22_X1 U61 ( .A1(A[8]), .A2(n67), .B1(B[8]), .B2(SEL), .ZN(n131) );
  INV_X1 U62 ( .A(n132), .ZN(Y[9]) );
  AOI22_X1 U63 ( .A1(A[9]), .A2(n67), .B1(SEL), .B2(B[9]), .ZN(n132) );
  INV_X1 U64 ( .A(n102), .ZN(Y[10]) );
  AOI22_X1 U65 ( .A1(A[10]), .A2(n33), .B1(B[10]), .B2(SEL), .ZN(n102) );
  INV_X1 U66 ( .A(n103), .ZN(Y[11]) );
  AOI22_X1 U67 ( .A1(A[11]), .A2(n33), .B1(B[11]), .B2(SEL), .ZN(n103) );
  INV_X1 U68 ( .A(SEL), .ZN(n100) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n33, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142;

  INV_X1 U1 ( .A(n111), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n122), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n68), .B1(B[1]), .B2(n74), .ZN(n122) );
  INV_X1 U4 ( .A(n141), .ZN(Y[8]) );
  INV_X1 U5 ( .A(n142), .ZN(Y[9]) );
  AOI22_X1 U6 ( .A1(A[9]), .A2(n68), .B1(n77), .B2(B[9]), .ZN(n142) );
  INV_X1 U7 ( .A(n139), .ZN(Y[6]) );
  AOI22_X1 U8 ( .A1(A[6]), .A2(n69), .B1(B[6]), .B2(n70), .ZN(n139) );
  INV_X1 U9 ( .A(n124), .ZN(Y[21]) );
  INV_X1 U10 ( .A(n133), .ZN(Y[2]) );
  AOI22_X1 U11 ( .A1(A[2]), .A2(n69), .B1(B[2]), .B2(n71), .ZN(n133) );
  INV_X1 U12 ( .A(n121), .ZN(Y[19]) );
  AOI22_X1 U13 ( .A1(A[19]), .A2(n68), .B1(B[19]), .B2(n75), .ZN(n121) );
  INV_X1 U14 ( .A(n132), .ZN(Y[29]) );
  AOI22_X1 U15 ( .A1(A[29]), .A2(n69), .B1(B[29]), .B2(n72), .ZN(n132) );
  INV_X1 U16 ( .A(n78), .ZN(n68) );
  INV_X1 U17 ( .A(n78), .ZN(n69) );
  INV_X1 U18 ( .A(n112), .ZN(Y[10]) );
  AOI22_X1 U19 ( .A1(A[10]), .A2(n68), .B1(B[10]), .B2(n77), .ZN(n112) );
  INV_X1 U20 ( .A(n136), .ZN(Y[3]) );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n68), .B1(B[3]), .B2(n71), .ZN(n136) );
  INV_X1 U22 ( .A(n129), .ZN(Y[26]) );
  AOI22_X1 U23 ( .A1(A[26]), .A2(n69), .B1(B[26]), .B2(n72), .ZN(n129) );
  INV_X1 U24 ( .A(n131), .ZN(Y[28]) );
  INV_X1 U25 ( .A(n137), .ZN(Y[4]) );
  AOI22_X1 U26 ( .A1(A[4]), .A2(n69), .B1(B[4]), .B2(n71), .ZN(n137) );
  INV_X1 U27 ( .A(n135), .ZN(Y[31]) );
  AOI22_X1 U28 ( .A1(A[31]), .A2(n68), .B1(B[31]), .B2(n71), .ZN(n135) );
  INV_X1 U29 ( .A(n113), .ZN(Y[11]) );
  AOI22_X1 U30 ( .A1(A[11]), .A2(n68), .B1(B[11]), .B2(n77), .ZN(n113) );
  INV_X1 U31 ( .A(n114), .ZN(Y[12]) );
  AOI22_X1 U32 ( .A1(A[12]), .A2(n68), .B1(B[12]), .B2(n76), .ZN(n114) );
  INV_X1 U33 ( .A(n115), .ZN(Y[13]) );
  INV_X1 U34 ( .A(n116), .ZN(Y[14]) );
  AOI22_X1 U35 ( .A1(A[14]), .A2(n68), .B1(B[14]), .B2(n76), .ZN(n116) );
  INV_X1 U36 ( .A(n117), .ZN(Y[15]) );
  AOI22_X1 U37 ( .A1(A[15]), .A2(n68), .B1(B[15]), .B2(n76), .ZN(n117) );
  INV_X1 U38 ( .A(n126), .ZN(Y[23]) );
  AOI22_X1 U39 ( .A1(A[23]), .A2(n69), .B1(B[23]), .B2(n73), .ZN(n126) );
  INV_X1 U40 ( .A(n119), .ZN(Y[17]) );
  AOI22_X1 U41 ( .A1(A[17]), .A2(n68), .B1(B[17]), .B2(n75), .ZN(n119) );
  INV_X1 U42 ( .A(n125), .ZN(Y[22]) );
  INV_X1 U43 ( .A(n118), .ZN(Y[16]) );
  AOI22_X1 U44 ( .A1(A[16]), .A2(n68), .B1(B[16]), .B2(n75), .ZN(n118) );
  INV_X1 U45 ( .A(n120), .ZN(Y[18]) );
  AOI22_X1 U46 ( .A1(A[18]), .A2(n68), .B1(B[18]), .B2(n75), .ZN(n120) );
  INV_X1 U47 ( .A(n138), .ZN(Y[5]) );
  AOI22_X1 U48 ( .A1(A[5]), .A2(n69), .B1(B[5]), .B2(n70), .ZN(n138) );
  INV_X1 U49 ( .A(n134), .ZN(Y[30]) );
  AOI22_X1 U50 ( .A1(A[30]), .A2(n69), .B1(B[30]), .B2(n74), .ZN(n134) );
  INV_X1 U51 ( .A(n130), .ZN(Y[27]) );
  AOI22_X1 U52 ( .A1(A[27]), .A2(n69), .B1(B[27]), .B2(n72), .ZN(n130) );
  INV_X1 U53 ( .A(n128), .ZN(Y[25]) );
  AOI22_X1 U54 ( .A1(A[25]), .A2(n69), .B1(B[25]), .B2(n73), .ZN(n128) );
  INV_X1 U55 ( .A(n123), .ZN(Y[20]) );
  AOI22_X1 U56 ( .A1(A[20]), .A2(n69), .B1(B[20]), .B2(n74), .ZN(n123) );
  INV_X1 U57 ( .A(n140), .ZN(Y[7]) );
  AOI22_X1 U58 ( .A1(A[7]), .A2(n68), .B1(B[7]), .B2(n70), .ZN(n140) );
  INV_X1 U59 ( .A(n127), .ZN(Y[24]) );
  AOI22_X1 U60 ( .A1(A[24]), .A2(n69), .B1(B[24]), .B2(n73), .ZN(n127) );
  BUF_X1 U61 ( .A(n66), .Z(n75) );
  BUF_X1 U62 ( .A(n33), .Z(n71) );
  BUF_X1 U63 ( .A(n67), .Z(n78) );
  BUF_X1 U64 ( .A(n33), .Z(n70) );
  BUF_X1 U65 ( .A(n67), .Z(n76) );
  BUF_X1 U66 ( .A(n66), .Z(n74) );
  BUF_X1 U67 ( .A(n33), .Z(n72) );
  BUF_X1 U68 ( .A(n66), .Z(n73) );
  BUF_X1 U69 ( .A(n67), .Z(n77) );
  BUF_X1 U70 ( .A(SEL), .Z(n66) );
  BUF_X1 U71 ( .A(SEL), .Z(n67) );
  BUF_X1 U72 ( .A(SEL), .Z(n33) );
  AOI22_X1 U73 ( .A1(A[13]), .A2(n68), .B1(B[13]), .B2(n76), .ZN(n115) );
  AOI22_X1 U74 ( .A1(A[22]), .A2(n69), .B1(B[22]), .B2(n73), .ZN(n125) );
  AOI22_X1 U75 ( .A1(A[28]), .A2(n69), .B1(B[28]), .B2(n72), .ZN(n131) );
  AOI22_X1 U76 ( .A1(A[21]), .A2(n69), .B1(B[21]), .B2(n74), .ZN(n124) );
  AOI22_X1 U77 ( .A1(A[0]), .A2(n68), .B1(B[0]), .B2(n77), .ZN(n111) );
  AOI22_X1 U78 ( .A1(A[8]), .A2(n69), .B1(B[8]), .B2(n70), .ZN(n141) );
endmodule


module PG_block_32 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_10 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module PG_block_31 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_30 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_29 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_28 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_27 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_26 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_25 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_24 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_23 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_22 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_21 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_20 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_19 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_18 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_17 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_16 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_15 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_14 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_13 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_12 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_11 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_10 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_9 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_8 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_7 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_6 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_5 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_4 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_3 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_2 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_1 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_9 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_27 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_8 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_26 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_25 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_24 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_23 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AOI21_X1 U1 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_22 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_21 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_20 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_19 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_18 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_17 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_16 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_15 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_14 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_13 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_12 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_11 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_10 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_9 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_8 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_7 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_6 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_G_7 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_5 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_6 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_5 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_4 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_3 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_2 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_1 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_4 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_3 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_2 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_1 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   Cin, first_generate, \p_vett[4][3] , \p_vett[4][2] , \p_vett[3][3] ,
         \p_vett[3][2] , \p_vett[3][1] , \p_vett[2][7] , \p_vett[2][6] ,
         \p_vett[2][5] , \p_vett[2][4] , \p_vett[2][3] , \p_vett[2][2] ,
         \p_vett[2][1] , \p_vett[1][15] , \p_vett[1][14] , \p_vett[1][13] ,
         \p_vett[1][12] , \p_vett[1][11] , \p_vett[1][10] , \p_vett[1][9] ,
         \p_vett[1][8] , \p_vett[1][7] , \p_vett[1][6] , \p_vett[1][5] ,
         \p_vett[1][4] , \p_vett[1][3] , \p_vett[1][2] , \p_vett[1][1] ,
         \p_vett[0][31] , \p_vett[0][30] , \p_vett[0][29] , \p_vett[0][28] ,
         \p_vett[0][27] , \p_vett[0][26] , \p_vett[0][25] , \p_vett[0][24] ,
         \p_vett[0][23] , \p_vett[0][22] , \p_vett[0][21] , \p_vett[0][20] ,
         \p_vett[0][19] , \p_vett[0][18] , \p_vett[0][17] , \p_vett[0][16] ,
         \p_vett[0][15] , \p_vett[0][14] , \p_vett[0][13] , \p_vett[0][12] ,
         \p_vett[0][11] , \p_vett[0][10] , \p_vett[0][9] , \p_vett[0][8] ,
         \p_vett[0][7] , \p_vett[0][6] , \p_vett[0][5] , \p_vett[0][4] ,
         \p_vett[0][3] , \p_vett[0][2] , \p_vett[0][1] , \p_vett[0][0] ,
         \g_vett[4][3] , \g_vett[4][2] , \g_vett[3][3] , \g_vett[3][2] ,
         \g_vett[3][1] , \g_vett[2][7] , \g_vett[2][6] , \g_vett[2][5] ,
         \g_vett[2][4] , \g_vett[2][3] , \g_vett[2][2] , \g_vett[2][1] ,
         \g_vett[1][15] , \g_vett[1][14] , \g_vett[1][13] , \g_vett[1][12] ,
         \g_vett[1][11] , \g_vett[1][10] , \g_vett[1][9] , \g_vett[1][8] ,
         \g_vett[1][7] , \g_vett[1][6] , \g_vett[1][5] , \g_vett[1][4] ,
         \g_vett[1][3] , \g_vett[1][2] , \g_vett[1][1] , \g_vett[1][0] ,
         \g_vett[0][31] , \g_vett[0][30] , \g_vett[0][29] , \g_vett[0][28] ,
         \g_vett[0][27] , \g_vett[0][26] , \g_vett[0][25] , \g_vett[0][24] ,
         \g_vett[0][23] , \g_vett[0][22] , \g_vett[0][21] , \g_vett[0][20] ,
         \g_vett[0][19] , \g_vett[0][18] , \g_vett[0][17] , \g_vett[0][16] ,
         \g_vett[0][15] , \g_vett[0][14] , \g_vett[0][13] , \g_vett[0][12] ,
         \g_vett[0][11] , \g_vett[0][10] , \g_vett[0][9] , \g_vett[0][8] ,
         \g_vett[0][7] , \g_vett[0][6] , \g_vett[0][5] , \g_vett[0][4] ,
         \g_vett[0][3] , \g_vett[0][2] , \g_vett[0][1] , \g_vett[0][0] ;
  assign Co[0] = Cin;

  PG_block_32 PGblock_first ( .A(A[0]), .B(B[0]), .G(first_generate), .P(
        \p_vett[0][0] ) );
  GENERAL_G_10 G_first ( .G_in(first_generate), .P_in(\p_vett[0][0] ), 
        .G_in_prev(Cin), .G_out(\g_vett[0][0] ) );
  PG_block_31 PG_0_1 ( .A(A[1]), .B(B[1]), .G(\g_vett[0][1] ), .P(
        \p_vett[0][1] ) );
  PG_block_30 PG_0_2 ( .A(A[2]), .B(B[2]), .G(\g_vett[0][2] ), .P(
        \p_vett[0][2] ) );
  PG_block_29 PG_0_3 ( .A(A[3]), .B(B[3]), .G(\g_vett[0][3] ), .P(
        \p_vett[0][3] ) );
  PG_block_28 PG_0_4 ( .A(A[4]), .B(B[4]), .G(\g_vett[0][4] ), .P(
        \p_vett[0][4] ) );
  PG_block_27 PG_0_5 ( .A(A[5]), .B(B[5]), .G(\g_vett[0][5] ), .P(
        \p_vett[0][5] ) );
  PG_block_26 PG_0_6 ( .A(A[6]), .B(B[6]), .G(\g_vett[0][6] ), .P(
        \p_vett[0][6] ) );
  PG_block_25 PG_0_7 ( .A(A[7]), .B(B[7]), .G(\g_vett[0][7] ), .P(
        \p_vett[0][7] ) );
  PG_block_24 PG_0_8 ( .A(A[8]), .B(B[8]), .G(\g_vett[0][8] ), .P(
        \p_vett[0][8] ) );
  PG_block_23 PG_0_9 ( .A(A[9]), .B(B[9]), .G(\g_vett[0][9] ), .P(
        \p_vett[0][9] ) );
  PG_block_22 PG_0_10 ( .A(A[10]), .B(B[10]), .G(\g_vett[0][10] ), .P(
        \p_vett[0][10] ) );
  PG_block_21 PG_0_11 ( .A(A[11]), .B(B[11]), .G(\g_vett[0][11] ), .P(
        \p_vett[0][11] ) );
  PG_block_20 PG_0_12 ( .A(A[12]), .B(B[12]), .G(\g_vett[0][12] ), .P(
        \p_vett[0][12] ) );
  PG_block_19 PG_0_13 ( .A(A[13]), .B(B[13]), .G(\g_vett[0][13] ), .P(
        \p_vett[0][13] ) );
  PG_block_18 PG_0_14 ( .A(A[14]), .B(B[14]), .G(\g_vett[0][14] ), .P(
        \p_vett[0][14] ) );
  PG_block_17 PG_0_15 ( .A(A[15]), .B(B[15]), .G(\g_vett[0][15] ), .P(
        \p_vett[0][15] ) );
  PG_block_16 PG_0_16 ( .A(A[16]), .B(B[16]), .G(\g_vett[0][16] ), .P(
        \p_vett[0][16] ) );
  PG_block_15 PG_0_17 ( .A(A[17]), .B(B[17]), .G(\g_vett[0][17] ), .P(
        \p_vett[0][17] ) );
  PG_block_14 PG_0_18 ( .A(A[18]), .B(B[18]), .G(\g_vett[0][18] ), .P(
        \p_vett[0][18] ) );
  PG_block_13 PG_0_19 ( .A(A[19]), .B(B[19]), .G(\g_vett[0][19] ), .P(
        \p_vett[0][19] ) );
  PG_block_12 PG_0_20 ( .A(A[20]), .B(B[20]), .G(\g_vett[0][20] ), .P(
        \p_vett[0][20] ) );
  PG_block_11 PG_0_21 ( .A(A[21]), .B(B[21]), .G(\g_vett[0][21] ), .P(
        \p_vett[0][21] ) );
  PG_block_10 PG_0_22 ( .A(A[22]), .B(B[22]), .G(\g_vett[0][22] ), .P(
        \p_vett[0][22] ) );
  PG_block_9 PG_0_23 ( .A(A[23]), .B(B[23]), .G(\g_vett[0][23] ), .P(
        \p_vett[0][23] ) );
  PG_block_8 PG_0_24 ( .A(A[24]), .B(B[24]), .G(\g_vett[0][24] ), .P(
        \p_vett[0][24] ) );
  PG_block_7 PG_0_25 ( .A(A[25]), .B(B[25]), .G(\g_vett[0][25] ), .P(
        \p_vett[0][25] ) );
  PG_block_6 PG_0_26 ( .A(A[26]), .B(B[26]), .G(\g_vett[0][26] ), .P(
        \p_vett[0][26] ) );
  PG_block_5 PG_0_27 ( .A(A[27]), .B(B[27]), .G(\g_vett[0][27] ), .P(
        \p_vett[0][27] ) );
  PG_block_4 PG_0_28 ( .A(A[28]), .B(B[28]), .G(\g_vett[0][28] ), .P(
        \p_vett[0][28] ) );
  PG_block_3 PG_0_29 ( .A(A[29]), .B(B[29]), .G(\g_vett[0][29] ), .P(
        \p_vett[0][29] ) );
  PG_block_2 PG_0_30 ( .A(A[30]), .B(B[30]), .G(\g_vett[0][30] ), .P(
        \p_vett[0][30] ) );
  PG_block_1 PG_0_31 ( .A(A[31]), .B(B[31]), .G(\g_vett[0][31] ), .P(
        \p_vett[0][31] ) );
  GENERAL_G_9 G_0_0_0 ( .G_in(\g_vett[0][1] ), .P_in(\p_vett[0][1] ), 
        .G_in_prev(\g_vett[0][0] ), .G_out(\g_vett[1][0] ) );
  GENERAL_PG_27 PG_1_0_0 ( .G_in(\g_vett[0][3] ), .P_in(\p_vett[0][3] ), 
        .G_in_prev(\g_vett[0][2] ), .P_in_prev(\p_vett[0][2] ), .G_out(
        \g_vett[1][1] ), .P_out(\p_vett[1][1] ) );
  GENERAL_G_8 G_1_0_0 ( .G_in(\g_vett[1][1] ), .P_in(\p_vett[1][1] ), 
        .G_in_prev(\g_vett[1][0] ), .G_out(Co[1]) );
  GENERAL_PG_26 PG_2_0_1 ( .G_in(\g_vett[0][5] ), .P_in(\p_vett[0][5] ), 
        .G_in_prev(\g_vett[0][4] ), .P_in_prev(\p_vett[0][4] ), .G_out(
        \g_vett[1][2] ), .P_out(\p_vett[1][2] ) );
  GENERAL_PG_25 PG_3_0_1 ( .G_in(\g_vett[0][7] ), .P_in(\p_vett[0][7] ), 
        .G_in_prev(\g_vett[0][6] ), .P_in_prev(\p_vett[0][6] ), .G_out(
        \g_vett[1][3] ), .P_out(\p_vett[1][3] ) );
  GENERAL_PG_24 PG_4_0_1 ( .G_in(\g_vett[1][3] ), .P_in(\p_vett[1][3] ), 
        .G_in_prev(\g_vett[1][2] ), .P_in_prev(\p_vett[1][2] ), .G_out(
        \g_vett[2][1] ), .P_out(\p_vett[2][1] ) );
  GENERAL_PG_23 PG_2_0_2 ( .G_in(\g_vett[0][9] ), .P_in(\p_vett[0][9] ), 
        .G_in_prev(\g_vett[0][8] ), .P_in_prev(\p_vett[0][8] ), .G_out(
        \g_vett[1][4] ), .P_out(\p_vett[1][4] ) );
  GENERAL_PG_22 PG_3_0_2 ( .G_in(\g_vett[0][11] ), .P_in(\p_vett[0][11] ), 
        .G_in_prev(\g_vett[0][10] ), .P_in_prev(\p_vett[0][10] ), .G_out(
        \g_vett[1][5] ), .P_out(\p_vett[1][5] ) );
  GENERAL_PG_21 PG_4_0_2 ( .G_in(\g_vett[1][5] ), .P_in(\p_vett[1][5] ), 
        .G_in_prev(\g_vett[1][4] ), .P_in_prev(\p_vett[1][4] ), .G_out(
        \g_vett[2][2] ), .P_out(\p_vett[2][2] ) );
  GENERAL_PG_20 PG_2_0_3 ( .G_in(\g_vett[0][13] ), .P_in(\p_vett[0][13] ), 
        .G_in_prev(\g_vett[0][12] ), .P_in_prev(\p_vett[0][12] ), .G_out(
        \g_vett[1][6] ), .P_out(\p_vett[1][6] ) );
  GENERAL_PG_19 PG_3_0_3 ( .G_in(\g_vett[0][15] ), .P_in(\p_vett[0][15] ), 
        .G_in_prev(\g_vett[0][14] ), .P_in_prev(\p_vett[0][14] ), .G_out(
        \g_vett[1][7] ), .P_out(\p_vett[1][7] ) );
  GENERAL_PG_18 PG_4_0_3 ( .G_in(\g_vett[1][7] ), .P_in(\p_vett[1][7] ), 
        .G_in_prev(\g_vett[1][6] ), .P_in_prev(\p_vett[1][6] ), .G_out(
        \g_vett[2][3] ), .P_out(\p_vett[2][3] ) );
  GENERAL_PG_17 PG_2_0_4 ( .G_in(\g_vett[0][17] ), .P_in(\p_vett[0][17] ), 
        .G_in_prev(\g_vett[0][16] ), .P_in_prev(\p_vett[0][16] ), .G_out(
        \g_vett[1][8] ), .P_out(\p_vett[1][8] ) );
  GENERAL_PG_16 PG_3_0_4 ( .G_in(\g_vett[0][19] ), .P_in(\p_vett[0][19] ), 
        .G_in_prev(\g_vett[0][18] ), .P_in_prev(\p_vett[0][18] ), .G_out(
        \g_vett[1][9] ), .P_out(\p_vett[1][9] ) );
  GENERAL_PG_15 PG_4_0_4 ( .G_in(\g_vett[1][9] ), .P_in(\p_vett[1][9] ), 
        .G_in_prev(\g_vett[1][8] ), .P_in_prev(\p_vett[1][8] ), .G_out(
        \g_vett[2][4] ), .P_out(\p_vett[2][4] ) );
  GENERAL_PG_14 PG_2_0_5 ( .G_in(\g_vett[0][21] ), .P_in(\p_vett[0][21] ), 
        .G_in_prev(\g_vett[0][20] ), .P_in_prev(\p_vett[0][20] ), .G_out(
        \g_vett[1][10] ), .P_out(\p_vett[1][10] ) );
  GENERAL_PG_13 PG_3_0_5 ( .G_in(\g_vett[0][23] ), .P_in(\p_vett[0][23] ), 
        .G_in_prev(\g_vett[0][22] ), .P_in_prev(\p_vett[0][22] ), .G_out(
        \g_vett[1][11] ), .P_out(\p_vett[1][11] ) );
  GENERAL_PG_12 PG_4_0_5 ( .G_in(\g_vett[1][11] ), .P_in(\p_vett[1][11] ), 
        .G_in_prev(\g_vett[1][10] ), .P_in_prev(\p_vett[1][10] ), .G_out(
        \g_vett[2][5] ), .P_out(\p_vett[2][5] ) );
  GENERAL_PG_11 PG_2_0_6 ( .G_in(\g_vett[0][25] ), .P_in(\p_vett[0][25] ), 
        .G_in_prev(\g_vett[0][24] ), .P_in_prev(\p_vett[0][24] ), .G_out(
        \g_vett[1][12] ), .P_out(\p_vett[1][12] ) );
  GENERAL_PG_10 PG_3_0_6 ( .G_in(\g_vett[0][27] ), .P_in(\p_vett[0][27] ), 
        .G_in_prev(\g_vett[0][26] ), .P_in_prev(\p_vett[0][26] ), .G_out(
        \g_vett[1][13] ), .P_out(\p_vett[1][13] ) );
  GENERAL_PG_9 PG_4_0_6 ( .G_in(\g_vett[1][13] ), .P_in(\p_vett[1][13] ), 
        .G_in_prev(\g_vett[1][12] ), .P_in_prev(\p_vett[1][12] ), .G_out(
        \g_vett[2][6] ), .P_out(\p_vett[2][6] ) );
  GENERAL_PG_8 PG_2_0_7 ( .G_in(\g_vett[0][29] ), .P_in(\p_vett[0][29] ), 
        .G_in_prev(\g_vett[0][28] ), .P_in_prev(\p_vett[0][28] ), .G_out(
        \g_vett[1][14] ), .P_out(\p_vett[1][14] ) );
  GENERAL_PG_7 PG_3_0_7 ( .G_in(\g_vett[0][31] ), .P_in(\p_vett[0][31] ), 
        .G_in_prev(\g_vett[0][30] ), .P_in_prev(\p_vett[0][30] ), .G_out(
        \g_vett[1][15] ), .P_out(\p_vett[1][15] ) );
  GENERAL_PG_6 PG_4_0_7 ( .G_in(\g_vett[1][15] ), .P_in(\p_vett[1][15] ), 
        .G_in_prev(\g_vett[1][14] ), .P_in_prev(\p_vett[1][14] ), .G_out(
        \g_vett[2][7] ), .P_out(\p_vett[2][7] ) );
  GENERAL_G_7 G_2_1_0 ( .G_in(\g_vett[2][1] ), .P_in(\p_vett[2][1] ), 
        .G_in_prev(Co[1]), .G_out(Co[2]) );
  GENERAL_PG_5 PG_5_1_0 ( .G_in(\g_vett[2][3] ), .P_in(\p_vett[2][3] ), 
        .G_in_prev(\g_vett[2][2] ), .P_in_prev(\p_vett[2][2] ), .G_out(
        \g_vett[3][1] ), .P_out(\p_vett[3][1] ) );
  GENERAL_G_6 G_3_1_0 ( .G_in(\g_vett[2][2] ), .P_in(\p_vett[2][2] ), 
        .G_in_prev(Co[2]), .G_out(Co[3]) );
  GENERAL_G_5 G_4_1_0 ( .G_in(\g_vett[3][1] ), .P_in(\p_vett[3][1] ), 
        .G_in_prev(Co[2]), .G_out(Co[4]) );
  GENERAL_PG_4 PG_6_1_1 ( .G_in(\g_vett[2][5] ), .P_in(\p_vett[2][5] ), 
        .G_in_prev(\g_vett[2][4] ), .P_in_prev(\p_vett[2][4] ), .G_out(
        \g_vett[3][2] ), .P_out(\p_vett[3][2] ) );
  GENERAL_PG_3 PG_7_1_1 ( .G_in(\g_vett[2][7] ), .P_in(\p_vett[2][7] ), 
        .G_in_prev(\g_vett[2][6] ), .P_in_prev(\p_vett[2][6] ), .G_out(
        \g_vett[3][3] ), .P_out(\p_vett[3][3] ) );
  GENERAL_PG_2 PG_8_1_1 ( .G_in(\g_vett[2][6] ), .P_in(\p_vett[2][6] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][2] ), .P_out(\p_vett[4][2] ) );
  GENERAL_PG_1 PG_9_1_1 ( .G_in(\g_vett[3][3] ), .P_in(\p_vett[3][3] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][3] ), .P_out(\p_vett[4][3] ) );
  GENERAL_G_4 G_5_2_0 ( .G_in(\g_vett[2][4] ), .P_in(\p_vett[2][4] ), 
        .G_in_prev(Co[4]), .G_out(Co[5]) );
  GENERAL_G_3 G_6_2_1 ( .G_in(\g_vett[3][2] ), .P_in(\p_vett[3][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[6]) );
  GENERAL_G_2 G_7_2_2 ( .G_in(\g_vett[4][2] ), .P_in(\p_vett[4][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[7]) );
  GENERAL_G_1 G_8_2_3 ( .G_in(\g_vett[4][3] ), .P_in(\p_vett[4][3] ), 
        .G_in_prev(Co[4]) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_16 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U2 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U5 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U7 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U9 ( .A(SEL), .ZN(n13) );
endmodule


module MUX21_GENERIC_NBIT4_15 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  INV_X1 U5 ( .A(SEL), .ZN(n13) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_8 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_16 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_15 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_16 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_15 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_14 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_13 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_7 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_14 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_13 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_14 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_13 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_12 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U4 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U6 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U8 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
endmodule


module MUX21_GENERIC_NBIT4_11 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_6 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_12 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_11 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_12 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_11 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_10 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U6 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U8 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
endmodule


module MUX21_GENERIC_NBIT4_9 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_5 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_10 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_9 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_10 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_9 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({1'b0, 
        1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_8 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U6 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_4 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_8 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_7 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_8 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_7 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({1'b0, 
        1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_3 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_6 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_5 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_6 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_5 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({1'b0, 
        1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U8 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_2 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_4 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_3 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_4 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_3 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({1'b0, 
        1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U8 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_1 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_2 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_1 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_2 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_1 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({1'b0, 
        1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module SUMGEN_NBIT32_NBLOCKS8_1 ( A, B, cin_vect, Co, SUM );
  input [31:0] A;
  input [31:0] B;
  input [7:0] cin_vect;
  output [31:0] SUM;
  output Co;


  CSblock_NBIT4_8 block_i_0 ( .A(A[3:0]), .B(B[3:0]), .cin(cin_vect[0]), .Y(
        SUM[3:0]) );
  CSblock_NBIT4_7 block_i_1 ( .A(A[7:4]), .B(B[7:4]), .cin(cin_vect[1]), .Y(
        SUM[7:4]) );
  CSblock_NBIT4_6 block_i_2 ( .A(A[11:8]), .B(B[11:8]), .cin(cin_vect[2]), .Y(
        SUM[11:8]) );
  CSblock_NBIT4_5 block_i_3 ( .A(A[15:12]), .B(B[15:12]), .cin(cin_vect[3]), 
        .Y(SUM[15:12]) );
  CSblock_NBIT4_4 block_i_4 ( .A(A[19:16]), .B(B[19:16]), .cin(cin_vect[4]), 
        .Y(SUM[19:16]) );
  CSblock_NBIT4_3 block_i_5 ( .A(A[23:20]), .B(B[23:20]), .cin(cin_vect[5]), 
        .Y(SUM[23:20]) );
  CSblock_NBIT4_2 block_i_6 ( .A(A[27:24]), .B(B[27:24]), .cin(cin_vect[6]), 
        .Y(SUM[27:24]) );
  CSblock_NBIT4_1 block_i_7 ( .A(A[31:28]), .B(B[31:28]), .cin(cin_vect[7]), 
        .Y(SUM[31:28]), .Co(Co) );
endmodule


module P4_ADDER_NBIT32_NBIT_PER_BLOCK4_1 ( A, B, Cin, Cout, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input Cin;
  output Cout;

  wire   [7:0] outCarryGen;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 CG ( .A(A), .B(B), .Cin(Cin), .Co(
        outCarryGen) );
  SUMGEN_NBIT32_NBLOCKS8_1 SG ( .A(A), .B(B), .cin_vect(outCarryGen), .Co(Cout), .SUM(Y) );
endmodule


module and_gate_nbit32 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;


  AND2_X1 U1 ( .A1(B[5]), .A2(A[5]), .ZN(Y[5]) );
  AND2_X1 U2 ( .A1(B[12]), .A2(A[12]), .ZN(Y[12]) );
  AND2_X1 U3 ( .A1(B[7]), .A2(A[7]), .ZN(Y[7]) );
  AND2_X1 U4 ( .A1(B[9]), .A2(A[9]), .ZN(Y[9]) );
  AND2_X1 U5 ( .A1(B[6]), .A2(A[6]), .ZN(Y[6]) );
  AND2_X1 U6 ( .A1(B[4]), .A2(A[4]), .ZN(Y[4]) );
  AND2_X1 U7 ( .A1(B[3]), .A2(A[3]), .ZN(Y[3]) );
  AND2_X1 U8 ( .A1(B[31]), .A2(A[31]), .ZN(Y[31]) );
  AND2_X1 U9 ( .A1(B[17]), .A2(A[17]), .ZN(Y[17]) );
  AND2_X1 U10 ( .A1(B[14]), .A2(A[14]), .ZN(Y[14]) );
  AND2_X1 U11 ( .A1(B[23]), .A2(A[23]), .ZN(Y[23]) );
  AND2_X1 U12 ( .A1(B[11]), .A2(A[11]), .ZN(Y[11]) );
  AND2_X1 U13 ( .A1(B[18]), .A2(A[18]), .ZN(Y[18]) );
  AND2_X1 U14 ( .A1(B[1]), .A2(A[1]), .ZN(Y[1]) );
  AND2_X1 U15 ( .A1(B[15]), .A2(A[15]), .ZN(Y[15]) );
  AND2_X1 U16 ( .A1(B[27]), .A2(A[27]), .ZN(Y[27]) );
  AND2_X1 U17 ( .A1(B[16]), .A2(A[16]), .ZN(Y[16]) );
  AND2_X1 U18 ( .A1(B[24]), .A2(A[24]), .ZN(Y[24]) );
  AND2_X1 U19 ( .A1(B[21]), .A2(A[21]), .ZN(Y[21]) );
  AND2_X1 U20 ( .A1(B[10]), .A2(A[10]), .ZN(Y[10]) );
  AND2_X1 U21 ( .A1(B[25]), .A2(A[25]), .ZN(Y[25]) );
  AND2_X1 U22 ( .A1(B[19]), .A2(A[19]), .ZN(Y[19]) );
  AND2_X1 U23 ( .A1(B[20]), .A2(A[20]), .ZN(Y[20]) );
  AND2_X1 U24 ( .A1(B[13]), .A2(A[13]), .ZN(Y[13]) );
  AND2_X1 U25 ( .A1(B[26]), .A2(A[26]), .ZN(Y[26]) );
  AND2_X1 U26 ( .A1(B[29]), .A2(A[29]), .ZN(Y[29]) );
  AND2_X1 U27 ( .A1(B[30]), .A2(A[30]), .ZN(Y[30]) );
  AND2_X1 U28 ( .A1(B[2]), .A2(A[2]), .ZN(Y[2]) );
  AND2_X1 U29 ( .A1(B[22]), .A2(A[22]), .ZN(Y[22]) );
  AND2_X1 U30 ( .A1(B[28]), .A2(A[28]), .ZN(Y[28]) );
  AND2_X1 U31 ( .A1(B[0]), .A2(A[0]), .ZN(Y[0]) );
  AND2_X1 U32 ( .A1(B[8]), .A2(A[8]), .ZN(Y[8]) );
endmodule


module or_gate_nbit32 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;


  OR2_X1 U1 ( .A1(A[31]), .A2(B[31]), .ZN(Y[31]) );
  OR2_X1 U2 ( .A1(A[6]), .A2(B[6]), .ZN(Y[6]) );
  OR2_X1 U3 ( .A1(A[4]), .A2(B[4]), .ZN(Y[4]) );
  OR2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(Y[7]) );
  OR2_X1 U5 ( .A1(A[9]), .A2(B[9]), .ZN(Y[9]) );
  OR2_X1 U6 ( .A1(A[5]), .A2(B[5]), .ZN(Y[5]) );
  OR2_X1 U7 ( .A1(A[3]), .A2(B[3]), .ZN(Y[3]) );
  OR2_X1 U8 ( .A1(A[30]), .A2(B[30]), .ZN(Y[30]) );
  OR2_X1 U9 ( .A1(A[21]), .A2(B[21]), .ZN(Y[21]) );
  OR2_X1 U10 ( .A1(A[20]), .A2(B[20]), .ZN(Y[20]) );
  OR2_X1 U11 ( .A1(A[29]), .A2(B[29]), .ZN(Y[29]) );
  OR2_X1 U12 ( .A1(A[25]), .A2(B[25]), .ZN(Y[25]) );
  OR2_X1 U13 ( .A1(A[26]), .A2(B[26]), .ZN(Y[26]) );
  OR2_X1 U14 ( .A1(A[27]), .A2(B[27]), .ZN(Y[27]) );
  OR2_X1 U15 ( .A1(A[23]), .A2(B[23]), .ZN(Y[23]) );
  OR2_X1 U16 ( .A1(A[24]), .A2(B[24]), .ZN(Y[24]) );
  OR2_X1 U17 ( .A1(A[15]), .A2(B[15]), .ZN(Y[15]) );
  OR2_X1 U18 ( .A1(A[10]), .A2(B[10]), .ZN(Y[10]) );
  OR2_X1 U19 ( .A1(A[13]), .A2(B[13]), .ZN(Y[13]) );
  OR2_X1 U20 ( .A1(A[14]), .A2(B[14]), .ZN(Y[14]) );
  OR2_X1 U21 ( .A1(A[11]), .A2(B[11]), .ZN(Y[11]) );
  OR2_X1 U22 ( .A1(A[16]), .A2(B[16]), .ZN(Y[16]) );
  OR2_X1 U23 ( .A1(A[12]), .A2(B[12]), .ZN(Y[12]) );
  OR2_X1 U24 ( .A1(A[17]), .A2(B[17]), .ZN(Y[17]) );
  OR2_X1 U25 ( .A1(A[18]), .A2(B[18]), .ZN(Y[18]) );
  OR2_X1 U26 ( .A1(A[19]), .A2(B[19]), .ZN(Y[19]) );
  OR2_X1 U27 ( .A1(A[1]), .A2(B[1]), .ZN(Y[1]) );
  OR2_X1 U28 ( .A1(A[2]), .A2(B[2]), .ZN(Y[2]) );
  OR2_X1 U29 ( .A1(A[22]), .A2(B[22]), .ZN(Y[22]) );
  OR2_X1 U30 ( .A1(A[28]), .A2(B[28]), .ZN(Y[28]) );
  OR2_X1 U31 ( .A1(A[0]), .A2(B[0]), .ZN(Y[0]) );
  OR2_X1 U32 ( .A1(A[8]), .A2(B[8]), .ZN(Y[8]) );
endmodule


module xor_gate_nbit32 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;


  XOR2_X1 U1 ( .A(B[9]), .B(A[9]), .Z(Y[9]) );
  XOR2_X1 U2 ( .A(B[8]), .B(A[8]), .Z(Y[8]) );
  XOR2_X1 U3 ( .A(B[7]), .B(A[7]), .Z(Y[7]) );
  XOR2_X1 U4 ( .A(B[6]), .B(A[6]), .Z(Y[6]) );
  XOR2_X1 U5 ( .A(B[5]), .B(A[5]), .Z(Y[5]) );
  XOR2_X1 U6 ( .A(B[4]), .B(A[4]), .Z(Y[4]) );
  XOR2_X1 U7 ( .A(B[3]), .B(A[3]), .Z(Y[3]) );
  XOR2_X1 U8 ( .A(B[31]), .B(A[31]), .Z(Y[31]) );
  XOR2_X1 U9 ( .A(B[30]), .B(A[30]), .Z(Y[30]) );
  XOR2_X1 U10 ( .A(B[2]), .B(A[2]), .Z(Y[2]) );
  XOR2_X1 U11 ( .A(B[29]), .B(A[29]), .Z(Y[29]) );
  XOR2_X1 U12 ( .A(B[28]), .B(A[28]), .Z(Y[28]) );
  XOR2_X1 U13 ( .A(B[27]), .B(A[27]), .Z(Y[27]) );
  XOR2_X1 U14 ( .A(B[26]), .B(A[26]), .Z(Y[26]) );
  XOR2_X1 U15 ( .A(B[25]), .B(A[25]), .Z(Y[25]) );
  XOR2_X1 U16 ( .A(B[24]), .B(A[24]), .Z(Y[24]) );
  XOR2_X1 U17 ( .A(B[23]), .B(A[23]), .Z(Y[23]) );
  XOR2_X1 U18 ( .A(B[22]), .B(A[22]), .Z(Y[22]) );
  XOR2_X1 U19 ( .A(B[21]), .B(A[21]), .Z(Y[21]) );
  XOR2_X1 U20 ( .A(B[20]), .B(A[20]), .Z(Y[20]) );
  XOR2_X1 U21 ( .A(B[1]), .B(A[1]), .Z(Y[1]) );
  XOR2_X1 U22 ( .A(B[19]), .B(A[19]), .Z(Y[19]) );
  XOR2_X1 U23 ( .A(B[18]), .B(A[18]), .Z(Y[18]) );
  XOR2_X1 U24 ( .A(B[17]), .B(A[17]), .Z(Y[17]) );
  XOR2_X1 U25 ( .A(B[16]), .B(A[16]), .Z(Y[16]) );
  XOR2_X1 U26 ( .A(B[15]), .B(A[15]), .Z(Y[15]) );
  XOR2_X1 U27 ( .A(B[14]), .B(A[14]), .Z(Y[14]) );
  XOR2_X1 U28 ( .A(B[13]), .B(A[13]), .Z(Y[13]) );
  XOR2_X1 U29 ( .A(B[12]), .B(A[12]), .Z(Y[12]) );
  XOR2_X1 U30 ( .A(B[11]), .B(A[11]), .Z(Y[11]) );
  XOR2_X1 U31 ( .A(B[10]), .B(A[10]), .Z(Y[10]) );
  XOR2_X1 U32 ( .A(B[0]), .B(A[0]), .Z(Y[0]) );
endmodule


module shifter_sx_nbit32 ( r1, r2, data_out );
  input [31:0] r1;
  input [31:0] r2;
  output [31:0] data_out;
  wire   N1155, N1156, N1157, N1158, N1159, N1160, N1162, N1163, N1164, N1165,
         N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175,
         N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n451, n452,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677;

  DLH_X1 \data_out_reg[31]  ( .G(1'b1), .D(n629), .Q(data_out[31]) );
  DLH_X1 \data_out_reg[30]  ( .G(1'b1), .D(N1185), .Q(data_out[30]) );
  DLH_X1 \data_out_reg[29]  ( .G(1'b1), .D(N1184), .Q(data_out[29]) );
  DLH_X1 \data_out_reg[28]  ( .G(1'b1), .D(N1183), .Q(data_out[28]) );
  DLH_X1 \data_out_reg[27]  ( .G(1'b1), .D(N1182), .Q(data_out[27]) );
  DLH_X1 \data_out_reg[26]  ( .G(1'b1), .D(N1181), .Q(data_out[26]) );
  DLH_X1 \data_out_reg[25]  ( .G(1'b1), .D(N1180), .Q(data_out[25]) );
  DLH_X1 \data_out_reg[24]  ( .G(1'b1), .D(N1179), .Q(data_out[24]) );
  DLH_X1 \data_out_reg[23]  ( .G(1'b1), .D(N1178), .Q(data_out[23]) );
  DLH_X1 \data_out_reg[22]  ( .G(1'b1), .D(N1177), .Q(data_out[22]) );
  DLH_X1 \data_out_reg[21]  ( .G(1'b1), .D(N1176), .Q(data_out[21]) );
  DLH_X1 \data_out_reg[20]  ( .G(1'b1), .D(N1175), .Q(data_out[20]) );
  DLH_X1 \data_out_reg[19]  ( .G(1'b1), .D(N1174), .Q(data_out[19]) );
  DLH_X1 \data_out_reg[18]  ( .G(1'b1), .D(N1173), .Q(data_out[18]) );
  DLH_X1 \data_out_reg[17]  ( .G(1'b1), .D(N1172), .Q(data_out[17]) );
  DLH_X1 \data_out_reg[16]  ( .G(1'b1), .D(N1171), .Q(data_out[16]) );
  DLH_X1 \data_out_reg[15]  ( .G(1'b1), .D(N1170), .Q(data_out[15]) );
  DLH_X1 \data_out_reg[14]  ( .G(1'b1), .D(N1169), .Q(data_out[14]) );
  DLH_X1 \data_out_reg[13]  ( .G(1'b1), .D(N1168), .Q(data_out[13]) );
  DLH_X1 \data_out_reg[12]  ( .G(1'b1), .D(N1167), .Q(data_out[12]) );
  DLH_X1 \data_out_reg[11]  ( .G(1'b1), .D(N1166), .Q(data_out[11]) );
  DLH_X1 \data_out_reg[10]  ( .G(1'b1), .D(N1165), .Q(data_out[10]) );
  DLH_X1 \data_out_reg[9]  ( .G(1'b1), .D(N1164), .Q(data_out[9]) );
  DLH_X1 \data_out_reg[8]  ( .G(1'b1), .D(N1163), .Q(data_out[8]) );
  DLH_X1 \data_out_reg[7]  ( .G(1'b1), .D(N1162), .Q(data_out[7]) );
  DLH_X1 \data_out_reg[6]  ( .G(1'b1), .D(n452), .Q(data_out[6]) );
  DLH_X1 \data_out_reg[5]  ( .G(1'b1), .D(N1160), .Q(data_out[5]) );
  DLH_X1 \data_out_reg[4]  ( .G(1'b1), .D(N1159), .Q(data_out[4]) );
  DLH_X1 \data_out_reg[3]  ( .G(1'b1), .D(N1158), .Q(data_out[3]) );
  DLH_X1 \data_out_reg[2]  ( .G(1'b1), .D(N1157), .Q(data_out[2]) );
  DLH_X1 \data_out_reg[1]  ( .G(1'b1), .D(N1156), .Q(data_out[1]) );
  DLH_X1 \data_out_reg[0]  ( .G(1'b1), .D(N1155), .Q(data_out[0]) );
  OR4_X2 U349 ( .A1(n87), .A2(n93), .A3(n664), .A4(n657), .ZN(n153) );
  NAND2_X2 U367 ( .A1(n440), .A2(n433), .ZN(n167) );
  OAI33_X1 U476 ( .A1(n557), .A2(n85), .A3(n86), .B1(n88), .B2(n87), .B3(n89), 
        .ZN(n84) );
  NAND3_X1 U477 ( .A1(n200), .A2(n201), .A3(n202), .ZN(n197) );
  NAND3_X1 U478 ( .A1(n354), .A2(n455), .A3(n485), .ZN(n353) );
  NAND3_X1 U480 ( .A1(n554), .A2(n515), .A3(n633), .ZN(n432) );
  NAND3_X1 U483 ( .A1(r2[0]), .A2(n469), .A3(r2[4]), .ZN(n86) );
  INV_X1 U3 ( .A(n667), .ZN(n455) );
  NAND3_X1 U4 ( .A1(n469), .A2(n672), .A3(r2[4]), .ZN(n168) );
  AOI221_X1 U5 ( .B1(n637), .B2(r1[24]), .C1(n638), .C2(r1[25]), .A(n209), 
        .ZN(n208) );
  NOR2_X1 U6 ( .A1(n671), .A2(r2[2]), .ZN(n437) );
  AOI221_X1 U7 ( .B1(r1[22]), .B2(n641), .C1(r1[23]), .C2(n457), .A(n210), 
        .ZN(n207) );
  AND2_X1 U8 ( .A1(n366), .A2(n530), .ZN(n471) );
  INV_X1 U9 ( .A(n355), .ZN(n653) );
  NAND2_X1 U10 ( .A1(n669), .A2(n433), .ZN(n355) );
  INV_X1 U11 ( .A(n286), .ZN(n659) );
  NAND3_X1 U12 ( .A1(n291), .A2(n161), .A3(n334), .ZN(n160) );
  BUF_X1 U13 ( .A(n107), .Z(n528) );
  OAI221_X1 U14 ( .B1(n548), .B2(n674), .C1(n539), .C2(n675), .A(n191), .ZN(
        n189) );
  OAI222_X1 U15 ( .A1(n673), .A2(n167), .B1(n168), .B2(n677), .C1(n676), .C2(
        n526), .ZN(n190) );
  NOR2_X1 U16 ( .A1(n670), .A2(r2[1]), .ZN(n442) );
  OAI222_X1 U17 ( .A1(n676), .A2(n167), .B1(n168), .B2(n611), .C1(n619), .C2(
        n526), .ZN(n166) );
  AOI221_X1 U18 ( .B1(n604), .B2(n666), .C1(n601), .C2(n659), .A(n147), .ZN(
        n136) );
  AOI221_X1 U19 ( .B1(n606), .B2(n666), .C1(n604), .C2(n659), .A(n115), .ZN(
        n96) );
  INV_X1 U20 ( .A(n471), .ZN(n129) );
  INV_X1 U21 ( .A(n466), .ZN(n363) );
  AOI221_X1 U22 ( .B1(n592), .B2(n653), .C1(r1[6]), .C2(n667), .A(n282), .ZN(
        n275) );
  AOI221_X1 U23 ( .B1(n586), .B2(n666), .C1(n581), .C2(n659), .A(n240), .ZN(
        n229) );
  AOI221_X1 U24 ( .B1(n590), .B2(n666), .C1(n586), .C2(n659), .A(n226), .ZN(
        n215) );
  AOI221_X1 U25 ( .B1(n592), .B2(n666), .C1(n590), .C2(n659), .A(n203), .ZN(
        n202) );
  INV_X1 U26 ( .A(n154), .ZN(n664) );
  OAI222_X1 U27 ( .A1(n569), .A2(n546), .B1(n431), .B2(n403), .C1(n576), .C2(
        n550), .ZN(N1158) );
  OAI221_X1 U28 ( .B1(n402), .B2(n403), .C1(n110), .C2(n557), .A(n404), .ZN(
        N1165) );
  AOI221_X1 U29 ( .B1(n636), .B2(n560), .C1(n648), .C2(n557), .A(n315), .ZN(
        n381) );
  AOI222_X1 U30 ( .A1(n648), .A2(n563), .B1(n359), .B2(n372), .C1(r1[2]), .C2(
        n636), .ZN(n371) );
  BUF_X1 U31 ( .A(n107), .Z(n529) );
  CLKBUF_X1 U32 ( .A(n128), .Z(n456) );
  AND2_X1 U33 ( .A1(n351), .A2(n642), .ZN(n457) );
  OR3_X1 U34 ( .A1(r2[5]), .A2(r2[31]), .A3(r2[30]), .ZN(n458) );
  AND2_X1 U35 ( .A1(n430), .A2(n471), .ZN(n459) );
  AND2_X1 U36 ( .A1(n103), .A2(n102), .ZN(n460) );
  OR3_X1 U37 ( .A1(r2[25]), .A2(r2[24]), .A3(r2[23]), .ZN(n461) );
  OR3_X1 U38 ( .A1(n188), .A2(n189), .A3(n190), .ZN(n462) );
  OR2_X1 U39 ( .A1(n518), .A2(n517), .ZN(n463) );
  OR2_X1 U40 ( .A1(n512), .A2(n511), .ZN(n464) );
  AND2_X1 U41 ( .A1(n111), .A2(n110), .ZN(n364) );
  AND4_X2 U42 ( .A1(n446), .A2(n467), .A3(n444), .A4(n445), .ZN(n439) );
  CLKBUF_X3 U43 ( .A(n174), .Z(n540) );
  CLKBUF_X1 U44 ( .A(n658), .Z(n465) );
  AND2_X1 U45 ( .A1(n113), .A2(n470), .ZN(n390) );
  BUF_X2 U46 ( .A(n434), .Z(n502) );
  AND2_X2 U47 ( .A1(n439), .A2(n468), .ZN(n434) );
  NAND2_X1 U48 ( .A1(n196), .A2(n654), .ZN(n315) );
  INV_X1 U49 ( .A(n86), .ZN(n661) );
  AND2_X2 U50 ( .A1(n437), .A2(n433), .ZN(n466) );
  NAND2_X1 U51 ( .A1(n661), .A2(n436), .ZN(n116) );
  NAND2_X1 U52 ( .A1(n661), .A2(n438), .ZN(n100) );
  NOR2_X1 U53 ( .A1(n448), .A2(n458), .ZN(n467) );
  AND2_X1 U54 ( .A1(n672), .A2(n668), .ZN(n468) );
  AND4_X2 U55 ( .A1(n447), .A2(n446), .A3(n444), .A4(n445), .ZN(n469) );
  AOI221_X1 U56 ( .B1(r1[22]), .B2(n637), .C1(r1[23]), .C2(n638), .A(n237), 
        .ZN(n236) );
  NOR2_X1 U57 ( .A1(n187), .A2(n462), .ZN(n185) );
  NAND2_X1 U58 ( .A1(n502), .A2(n436), .ZN(n366) );
  OR2_X1 U59 ( .A1(n627), .A2(n494), .ZN(n509) );
  AND3_X1 U60 ( .A1(n283), .A2(n355), .A3(n168), .ZN(n470) );
  AND2_X1 U61 ( .A1(n524), .A2(n167), .ZN(n443) );
  INV_X1 U62 ( .A(n167), .ZN(n650) );
  INV_X1 U63 ( .A(n111), .ZN(n652) );
  NAND2_X1 U64 ( .A1(n632), .A2(n459), .ZN(n429) );
  NAND2_X1 U65 ( .A1(n666), .A2(r2[3]), .ZN(n472) );
  AND3_X2 U66 ( .A1(n390), .A2(n364), .A3(n527), .ZN(n351) );
  NAND2_X2 U67 ( .A1(n435), .A2(n502), .ZN(n110) );
  AND3_X1 U68 ( .A1(n364), .A2(n390), .A3(n527), .ZN(n473) );
  AND3_X1 U69 ( .A1(n364), .A2(n390), .A3(n527), .ZN(n500) );
  OR2_X1 U70 ( .A1(n627), .A2(n544), .ZN(n474) );
  OR2_X1 U71 ( .A1(n628), .A2(n550), .ZN(n475) );
  NAND3_X1 U72 ( .A1(n474), .A2(n475), .A3(n130), .ZN(N1185) );
  CLKBUF_X1 U73 ( .A(n640), .Z(n476) );
  INV_X1 U74 ( .A(n528), .ZN(n640) );
  AND2_X1 U75 ( .A1(n551), .A2(n657), .ZN(n477) );
  AND2_X1 U76 ( .A1(n664), .A2(n561), .ZN(n478) );
  NOR3_X1 U77 ( .A1(n477), .A2(n478), .A3(n228), .ZN(n227) );
  NAND2_X1 U78 ( .A1(n654), .A2(n231), .ZN(n479) );
  NAND2_X1 U79 ( .A1(n590), .A2(n655), .ZN(n480) );
  INV_X1 U80 ( .A(n232), .ZN(n481) );
  AND3_X1 U81 ( .A1(n479), .A2(n480), .A3(n481), .ZN(n230) );
  INV_X1 U82 ( .A(n199), .ZN(n657) );
  OR2_X1 U83 ( .A1(n84), .A2(n464), .ZN(n629) );
  NAND2_X1 U84 ( .A1(r1[26]), .A2(n641), .ZN(n482) );
  NAND2_X1 U85 ( .A1(r1[27]), .A2(n457), .ZN(n483) );
  INV_X1 U86 ( .A(n109), .ZN(n484) );
  AND3_X1 U87 ( .A1(n482), .A2(n483), .A3(n484), .ZN(n104) );
  CLKBUF_X1 U88 ( .A(n634), .Z(n485) );
  CLKBUF_X1 U89 ( .A(n93), .Z(n486) );
  OR2_X1 U90 ( .A1(n588), .A2(n546), .ZN(n487) );
  OR2_X1 U91 ( .A1(n591), .A2(n550), .ZN(n488) );
  NAND3_X1 U92 ( .A1(n487), .A2(n488), .A3(n123), .ZN(n452) );
  AOI221_X1 U93 ( .B1(r1[16]), .B2(n641), .C1(r1[17]), .C2(n457), .A(n298), 
        .ZN(n295) );
  AOI221_X1 U94 ( .B1(r1[20]), .B2(n641), .C1(n618), .C2(n457), .A(n238), .ZN(
        n235) );
  AOI221_X1 U95 ( .B1(n617), .B2(n641), .C1(r1[22]), .C2(n457), .A(n224), .ZN(
        n221) );
  NOR3_X1 U96 ( .A1(r2[11]), .A2(r2[12]), .A3(r2[10]), .ZN(n489) );
  NOR2_X1 U97 ( .A1(n451), .A2(n490), .ZN(n444) );
  INV_X1 U98 ( .A(n489), .ZN(n490) );
  AND2_X1 U99 ( .A1(n491), .A2(n522), .ZN(n445) );
  NOR4_X1 U100 ( .A1(r2[20]), .A2(r2[19]), .A3(r2[22]), .A4(r2[21]), .ZN(n491)
         );
  OR2_X1 U101 ( .A1(n623), .A2(n540), .ZN(n492) );
  OR2_X1 U102 ( .A1(n538), .A2(n624), .ZN(n493) );
  NAND3_X1 U103 ( .A1(n193), .A2(n493), .A3(n492), .ZN(n187) );
  BUF_X2 U104 ( .A(n175), .Z(n538) );
  NAND2_X1 U105 ( .A1(n515), .A2(n351), .ZN(n494) );
  NOR2_X2 U106 ( .A1(n153), .A2(n89), .ZN(n196) );
  OR2_X1 U107 ( .A1(n676), .A2(n545), .ZN(n495) );
  OR2_X1 U108 ( .A1(n619), .A2(n550), .ZN(n496) );
  NAND3_X1 U109 ( .A1(n495), .A2(n496), .A3(n284), .ZN(N1176) );
  NAND2_X1 U110 ( .A1(n579), .A2(n656), .ZN(n497) );
  NAND2_X1 U111 ( .A1(n291), .A2(n292), .ZN(n498) );
  NAND2_X1 U112 ( .A1(n571), .A2(n663), .ZN(n499) );
  AND3_X1 U113 ( .A1(n497), .A2(n498), .A3(n499), .ZN(n290) );
  INV_X1 U114 ( .A(n100), .ZN(n656) );
  AND2_X1 U115 ( .A1(n521), .A2(n520), .ZN(n501) );
  AND2_X1 U116 ( .A1(n519), .A2(n501), .ZN(n97) );
  NOR2_X1 U117 ( .A1(n95), .A2(n463), .ZN(n92) );
  INV_X1 U118 ( .A(n110), .ZN(n645) );
  OAI221_X4 U119 ( .B1(n111), .B2(n577), .C1(n110), .C2(n585), .A(n373), .ZN(
        n372) );
  AND2_X1 U120 ( .A1(n586), .A2(n657), .ZN(n503) );
  AND2_X1 U121 ( .A1(n590), .A2(n664), .ZN(n504) );
  NOR3_X1 U122 ( .A1(n135), .A2(n504), .A3(n503), .ZN(n133) );
  AND2_X1 U123 ( .A1(r1[27]), .A2(n637), .ZN(n505) );
  AND2_X1 U124 ( .A1(n638), .A2(r1[28]), .ZN(n506) );
  NOR3_X1 U125 ( .A1(n505), .A2(n506), .A3(n144), .ZN(n143) );
  NAND2_X1 U126 ( .A1(n667), .A2(n436), .ZN(n117) );
  INV_X2 U127 ( .A(n283), .ZN(n507) );
  NAND2_X1 U128 ( .A1(r1[28]), .A2(n637), .ZN(n508) );
  INV_X1 U129 ( .A(n106), .ZN(n510) );
  AND3_X1 U130 ( .A1(n508), .A2(n510), .A3(n509), .ZN(n105) );
  AND2_X1 U131 ( .A1(r1[30]), .A2(n646), .ZN(n511) );
  AND2_X1 U132 ( .A1(r1[31]), .A2(n523), .ZN(n512) );
  NOR2_X1 U133 ( .A1(n448), .A2(n458), .ZN(n447) );
  CLKBUF_X1 U134 ( .A(n364), .Z(n513) );
  INV_X1 U135 ( .A(n124), .ZN(n514) );
  NAND3_X1 U136 ( .A1(n105), .A2(n104), .A3(n460), .ZN(n98) );
  INV_X1 U137 ( .A(n531), .ZN(n649) );
  OR4_X2 U138 ( .A1(r2[7]), .A2(r2[6]), .A3(r2[8]), .A4(r2[9]), .ZN(n448) );
  NAND2_X1 U139 ( .A1(n666), .A2(r2[3]), .ZN(n120) );
  AND2_X1 U140 ( .A1(n437), .A2(r2[3]), .ZN(n435) );
  AND4_X2 U141 ( .A1(n128), .A2(n471), .A3(n443), .A4(n417), .ZN(n515) );
  AND2_X1 U142 ( .A1(r2[0]), .A2(n668), .ZN(n516) );
  AND2_X2 U143 ( .A1(n439), .A2(n516), .ZN(n433) );
  AND2_X1 U144 ( .A1(n590), .A2(n657), .ZN(n517) );
  AND2_X1 U145 ( .A1(n592), .A2(n664), .ZN(n518) );
  NAND2_X1 U146 ( .A1(n98), .A2(n654), .ZN(n519) );
  NAND2_X1 U147 ( .A1(n542), .A2(n655), .ZN(n520) );
  INV_X1 U148 ( .A(n99), .ZN(n521) );
  NOR3_X1 U149 ( .A1(r2[17]), .A2(r2[18]), .A3(r2[16]), .ZN(n522) );
  INV_X2 U150 ( .A(n289), .ZN(n666) );
  INV_X2 U151 ( .A(n367), .ZN(n642) );
  INV_X2 U152 ( .A(n101), .ZN(n663) );
  NOR2_X2 U153 ( .A1(n670), .A2(n671), .ZN(n436) );
  CLKBUF_X1 U154 ( .A(n114), .Z(n547) );
  CLKBUF_X1 U155 ( .A(r1[0]), .Z(n555) );
  CLKBUF_X1 U156 ( .A(r1[0]), .Z(n556) );
  NOR2_X1 U157 ( .A1(n449), .A2(n461), .ZN(n446) );
  INV_X1 U158 ( .A(n160), .ZN(n654) );
  INV_X1 U159 ( .A(n315), .ZN(n634) );
  INV_X1 U160 ( .A(n161), .ZN(n655) );
  INV_X1 U161 ( .A(n534), .ZN(n639) );
  NOR2_X1 U162 ( .A1(n663), .A2(n656), .ZN(n291) );
  INV_X1 U163 ( .A(n196), .ZN(n631) );
  NAND2_X1 U164 ( .A1(n196), .A2(n334), .ZN(n270) );
  NOR2_X1 U165 ( .A1(n557), .A2(n550), .ZN(N1155) );
  INV_X1 U166 ( .A(n366), .ZN(n643) );
  INV_X1 U167 ( .A(n117), .ZN(n662) );
  INV_X1 U168 ( .A(n426), .ZN(n632) );
  AND4_X1 U169 ( .A1(n117), .A2(n116), .A3(n289), .A4(n286), .ZN(n334) );
  INV_X1 U170 ( .A(n121), .ZN(n646) );
  NAND2_X1 U171 ( .A1(n437), .A2(n661), .ZN(n161) );
  NAND2_X1 U172 ( .A1(n437), .A2(n667), .ZN(n101) );
  OAI22_X1 U173 ( .A1(n100), .A2(n614), .B1(n101), .B2(n611), .ZN(n99) );
  AOI22_X1 U174 ( .A1(n573), .A2(n666), .B1(r1[2]), .B2(n659), .ZN(n258) );
  AOI22_X1 U175 ( .A1(n581), .A2(n666), .B1(n573), .B2(n659), .ZN(n245) );
  INV_X1 U176 ( .A(n554), .ZN(n557) );
  AOI22_X1 U177 ( .A1(n580), .A2(n657), .B1(n553), .B2(n465), .ZN(n155) );
  AOI22_X1 U178 ( .A1(n573), .A2(n657), .B1(n665), .B2(n565), .ZN(n181) );
  AOI22_X1 U179 ( .A1(n573), .A2(n665), .B1(n660), .B2(n565), .ZN(n151) );
  OAI22_X1 U180 ( .A1(n560), .A2(n550), .B1(n557), .B2(n543), .ZN(N1156) );
  NAND2_X1 U181 ( .A1(n442), .A2(n667), .ZN(n289) );
  NAND2_X1 U182 ( .A1(n442), .A2(n661), .ZN(n286) );
  INV_X1 U183 ( .A(n582), .ZN(n585) );
  NAND2_X1 U184 ( .A1(n442), .A2(n434), .ZN(n367) );
  INV_X1 U185 ( .A(n119), .ZN(n665) );
  NAND2_X1 U186 ( .A1(n667), .A2(n669), .ZN(n94) );
  NAND2_X1 U187 ( .A1(n434), .A2(n669), .ZN(n283) );
  INV_X1 U188 ( .A(n403), .ZN(n633) );
  CLKBUF_X1 U189 ( .A(n172), .Z(n532) );
  BUF_X1 U190 ( .A(n121), .Z(n543) );
  CLKBUF_X1 U191 ( .A(n121), .Z(n544) );
  CLKBUF_X1 U192 ( .A(n108), .Z(n535) );
  CLKBUF_X1 U193 ( .A(n172), .Z(n533) );
  CLKBUF_X1 U194 ( .A(n121), .Z(n545) );
  CLKBUF_X1 U195 ( .A(n121), .Z(n546) );
  INV_X1 U196 ( .A(n118), .ZN(n660) );
  INV_X1 U197 ( .A(n564), .ZN(n560) );
  AOI211_X1 U198 ( .C1(n137), .C2(n136), .A(n657), .B(n664), .ZN(n135) );
  AOI22_X1 U199 ( .A1(n590), .A2(n652), .B1(n592), .B2(n645), .ZN(n342) );
  AOI22_X1 U200 ( .A1(n592), .A2(n652), .B1(n597), .B2(n645), .ZN(n332) );
  OAI222_X1 U201 ( .A1(n118), .A2(n578), .B1(n119), .B2(n585), .C1(n569), .C2(
        n472), .ZN(n132) );
  AOI221_X1 U202 ( .B1(n592), .B2(n507), .C1(r1[6]), .C2(n653), .A(n299), .ZN(
        n294) );
  AOI221_X1 U203 ( .B1(n606), .B2(n507), .C1(n604), .C2(n653), .A(n239), .ZN(
        n234) );
  INV_X1 U204 ( .A(n613), .ZN(n614) );
  OAI221_X1 U205 ( .B1(n324), .B2(n270), .C1(n325), .C2(n315), .A(n326), .ZN(
        N1173) );
  AOI22_X1 U206 ( .A1(n646), .A2(r1[17]), .B1(n523), .B2(r1[18]), .ZN(n326) );
  AOI22_X1 U207 ( .A1(n552), .A2(n663), .B1(n656), .B2(n562), .ZN(n324) );
  NOR4_X1 U208 ( .A1(n327), .A2(n328), .A3(n329), .A4(n330), .ZN(n325) );
  INV_X1 U209 ( .A(n601), .ZN(n603) );
  AOI22_X1 U210 ( .A1(n515), .A2(n561), .B1(n553), .B2(n466), .ZN(n431) );
  OAI221_X1 U211 ( .B1(n540), .B2(n619), .C1(n538), .C2(n620), .A(n254), .ZN(
        n248) );
  AOI22_X1 U212 ( .A1(r1[17]), .A2(n639), .B1(r1[18]), .B2(n640), .ZN(n254) );
  OAI221_X1 U213 ( .B1(n540), .B2(n611), .C1(n538), .C2(n614), .A(n352), .ZN(
        n345) );
  AOI22_X1 U214 ( .A1(n600), .A2(n639), .B1(n604), .B2(n476), .ZN(n352) );
  INV_X1 U215 ( .A(n610), .ZN(n611) );
  OAI22_X1 U216 ( .A1(n116), .A2(n568), .B1(n117), .B2(n576), .ZN(n240) );
  OAI22_X1 U217 ( .A1(n116), .A2(n575), .B1(n117), .B2(n585), .ZN(n226) );
  OAI221_X1 U218 ( .B1(n268), .B2(n631), .C1(n269), .C2(n270), .A(n271), .ZN(
        N1177) );
  AOI22_X1 U219 ( .A1(n646), .A2(n617), .B1(n523), .B2(r1[22]), .ZN(n271) );
  AOI222_X1 U220 ( .A1(n551), .A2(n662), .B1(n565), .B2(n666), .C1(n659), .C2(
        n563), .ZN(n268) );
  AOI221_X1 U221 ( .B1(n579), .B2(n663), .C1(n573), .C2(n655), .A(n272), .ZN(
        n269) );
  OAI221_X1 U222 ( .B1(n560), .B2(n545), .C1(n570), .C2(n550), .A(n432), .ZN(
        N1157) );
  OAI221_X1 U223 ( .B1(n575), .B2(n545), .C1(n585), .C2(n550), .A(n429), .ZN(
        N1159) );
  OAI221_X1 U224 ( .B1(n677), .B2(n544), .C1(n611), .C2(n550), .A(n379), .ZN(
        N1168) );
  NAND4_X1 U225 ( .A1(n355), .A2(n455), .A3(n380), .A4(n381), .ZN(n379) );
  AOI21_X1 U226 ( .B1(n359), .B2(n382), .A(n507), .ZN(n380) );
  OAI221_X1 U227 ( .B1(n611), .B2(n545), .C1(n614), .C2(n550), .A(n369), .ZN(
        N1169) );
  NAND4_X1 U228 ( .A1(n485), .A2(n370), .A3(n355), .A4(n455), .ZN(n369) );
  OAI22_X1 U229 ( .A1(n283), .A2(n557), .B1(n507), .B2(n371), .ZN(n370) );
  OAI21_X1 U230 ( .B1(n85), .B2(n86), .A(n543), .ZN(n87) );
  NAND2_X1 U231 ( .A1(n435), .A2(n661), .ZN(n118) );
  AOI22_X1 U232 ( .A1(n586), .A2(n663), .B1(r1[6]), .B2(n656), .ZN(n260) );
  INV_X1 U233 ( .A(n578), .ZN(n573) );
  INV_X1 U234 ( .A(n568), .ZN(n565) );
  NAND2_X1 U235 ( .A1(n435), .A2(n667), .ZN(n119) );
  INV_X1 U236 ( .A(n598), .ZN(n599) );
  NAND2_X1 U237 ( .A1(n440), .A2(n667), .ZN(n154) );
  AOI21_X1 U238 ( .B1(n636), .B2(n574), .A(n507), .ZN(n358) );
  AOI22_X1 U239 ( .A1(r1[17]), .A2(n652), .B1(r1[18]), .B2(n645), .ZN(n192) );
  NAND4_X1 U240 ( .A1(n120), .A2(n94), .A3(n118), .A4(n441), .ZN(n93) );
  NOR2_X1 U241 ( .A1(n665), .A2(n658), .ZN(n441) );
  AOI22_X1 U242 ( .A1(n581), .A2(n667), .B1(n606), .B2(n650), .ZN(n309) );
  AOI22_X1 U243 ( .A1(n600), .A2(n507), .B1(n597), .B2(n653), .ZN(n265) );
  AOI22_X1 U244 ( .A1(n590), .A2(n507), .B1(n586), .B2(n653), .ZN(n310) );
  AOI22_X1 U245 ( .A1(n612), .A2(n507), .B1(n610), .B2(n653), .ZN(n191) );
  AOI22_X1 U246 ( .A1(n565), .A2(n507), .B1(n653), .B2(n562), .ZN(n349) );
  OAI211_X1 U247 ( .C1(n363), .C2(n585), .A(n471), .B(n424), .ZN(n423) );
  INV_X1 U248 ( .A(r2[1]), .ZN(n671) );
  AND2_X1 U249 ( .A1(n434), .A2(n438), .ZN(n523) );
  INV_X1 U250 ( .A(r2[2]), .ZN(n670) );
  INV_X1 U251 ( .A(n85), .ZN(n669) );
  BUF_X1 U252 ( .A(n556), .Z(n551) );
  BUF_X1 U253 ( .A(n583), .Z(n581) );
  INV_X1 U254 ( .A(n134), .ZN(n658) );
  NAND2_X1 U255 ( .A1(n440), .A2(n661), .ZN(n199) );
  BUF_X1 U256 ( .A(n555), .Z(n553) );
  BUF_X1 U257 ( .A(n584), .Z(n580) );
  BUF_X1 U258 ( .A(n584), .Z(n579) );
  BUF_X1 U259 ( .A(n556), .Z(n552) );
  BUF_X1 U260 ( .A(n555), .Z(n554) );
  BUF_X1 U261 ( .A(n583), .Z(n582) );
  AOI221_X1 U262 ( .B1(n592), .B2(n649), .C1(n596), .C2(n642), .A(n395), .ZN(
        n391) );
  OAI22_X1 U263 ( .A1(n528), .A2(n673), .B1(n535), .B2(n616), .ZN(n237) );
  AOI22_X1 U264 ( .A1(n560), .A2(n651), .B1(n417), .B2(n418), .ZN(n416) );
  INV_X1 U265 ( .A(n605), .ZN(n604) );
  NOR3_X1 U266 ( .A1(r2[2]), .A2(r2[3]), .A3(r2[1]), .ZN(n438) );
  INV_X1 U267 ( .A(n587), .ZN(n586) );
  OAI221_X1 U268 ( .B1(n366), .B2(n603), .C1(n367), .C2(n607), .A(n368), .ZN(
        n361) );
  AOI22_X1 U269 ( .A1(n608), .A2(n652), .B1(n613), .B2(n645), .ZN(n253) );
  AOI22_X1 U270 ( .A1(n600), .A2(n652), .B1(n604), .B2(n645), .ZN(n311) );
  INV_X1 U271 ( .A(n607), .ZN(n606) );
  AOI22_X1 U272 ( .A1(n586), .A2(n652), .B1(r1[6]), .B2(n645), .ZN(n350) );
  AOI22_X1 U273 ( .A1(n596), .A2(n652), .B1(n602), .B2(n645), .ZN(n322) );
  INV_X1 U274 ( .A(n594), .ZN(n592) );
  NOR4_X1 U275 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(n259) );
  OAI221_X1 U276 ( .B1(n547), .B2(n607), .C1(n539), .C2(n605), .A(n265), .ZN(
        n263) );
  NOR4_X1 U277 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(n159) );
  OAI221_X1 U278 ( .B1(n547), .B2(n615), .C1(n539), .C2(n674), .A(n170), .ZN(
        n165) );
  OAI222_X1 U279 ( .A1(n585), .A2(n545), .B1(n425), .B2(n426), .C1(n588), .C2(
        n550), .ZN(N1160) );
  AOI22_X1 U280 ( .A1(n456), .A2(n574), .B1(n466), .B2(n567), .ZN(n428) );
  OAI222_X1 U281 ( .A1(n605), .A2(n544), .B1(n396), .B2(n397), .C1(n607), .C2(
        n550), .ZN(N1166) );
  OAI22_X1 U282 ( .A1(n116), .A2(n599), .B1(n117), .B2(n603), .ZN(n115) );
  OAI222_X1 U283 ( .A1(n675), .A2(n543), .B1(n344), .B2(n315), .C1(n674), .C2(
        n550), .ZN(N1171) );
  NOR4_X1 U284 ( .A1(n345), .A2(n346), .A3(n347), .A4(n348), .ZN(n344) );
  OAI221_X1 U285 ( .B1(n548), .B2(n585), .C1(n539), .C2(n577), .A(n349), .ZN(
        n347) );
  AOI221_X1 U286 ( .B1(n586), .B2(n651), .C1(r1[6]), .C2(n643), .A(n394), .ZN(
        n392) );
  AOI221_X1 U287 ( .B1(n656), .B2(n577), .C1(n663), .C2(n566), .A(n304), .ZN(
        n303) );
  NOR4_X1 U288 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n304) );
  OAI221_X1 U289 ( .B1(n114), .B2(n599), .C1(n539), .C2(n593), .A(n310), .ZN(
        n307) );
  AOI221_X1 U290 ( .B1(n542), .B2(n507), .C1(n606), .C2(n653), .A(n225), .ZN(
        n220) );
  INV_X1 U291 ( .A(n591), .ZN(n590) );
  OAI222_X1 U292 ( .A1(n118), .A2(n585), .B1(n119), .B2(n589), .C1(n472), .C2(
        n574), .ZN(n90) );
  OAI221_X1 U293 ( .B1(n246), .B2(n160), .C1(n161), .C2(n588), .A(n247), .ZN(
        n243) );
  AOI22_X1 U294 ( .A1(n590), .A2(n663), .B1(n592), .B2(n656), .ZN(n247) );
  NOR4_X1 U295 ( .A1(n248), .A2(n249), .A3(n250), .A4(n251), .ZN(n246) );
  OAI222_X1 U296 ( .A1(n675), .A2(n167), .B1(n455), .B2(n599), .C1(n674), .C2(
        n525), .ZN(n251) );
  OAI221_X1 U297 ( .B1(n540), .B2(n615), .C1(n538), .C2(n616), .A(n312), .ZN(
        n305) );
  AOI22_X1 U298 ( .A1(n608), .A2(n639), .B1(n613), .B2(n640), .ZN(n312) );
  OAI221_X1 U299 ( .B1(n540), .B2(n624), .C1(n538), .C2(n625), .A(n176), .ZN(
        n163) );
  AOI22_X1 U300 ( .A1(r1[22]), .A2(n639), .B1(r1[23]), .B2(n640), .ZN(n176) );
  OAI221_X1 U301 ( .B1(n540), .B2(n614), .C1(n538), .C2(n675), .A(n343), .ZN(
        n337) );
  AOI22_X1 U302 ( .A1(n604), .A2(n639), .B1(n606), .B2(n476), .ZN(n343) );
  OAI221_X1 U303 ( .B1(n540), .B2(n675), .C1(n538), .C2(n674), .A(n333), .ZN(
        n327) );
  AOI22_X1 U304 ( .A1(n606), .A2(n639), .B1(n542), .B2(n476), .ZN(n333) );
  OAI221_X1 U305 ( .B1(n540), .B2(n674), .C1(n538), .C2(n615), .A(n323), .ZN(
        n317) );
  AOI22_X1 U306 ( .A1(n542), .A2(n639), .B1(n609), .B2(n476), .ZN(n323) );
  AOI22_X1 U307 ( .A1(n617), .A2(n639), .B1(r1[22]), .B2(n640), .ZN(n193) );
  INV_X1 U308 ( .A(n542), .ZN(n677) );
  OAI22_X1 U309 ( .A1(n116), .A2(n593), .B1(n117), .B2(n599), .ZN(n147) );
  OAI22_X1 U310 ( .A1(n116), .A2(n585), .B1(n117), .B2(n587), .ZN(n203) );
  OAI221_X1 U311 ( .B1(n366), .B2(n589), .C1(n367), .C2(n594), .A(n401), .ZN(
        n398) );
  OAI221_X1 U312 ( .B1(n366), .B2(n595), .C1(n367), .C2(n603), .A(n386), .ZN(
        n383) );
  OAI221_X1 U313 ( .B1(n673), .B2(n543), .C1(n676), .C2(n550), .A(n300), .ZN(
        N1175) );
  NAND4_X1 U314 ( .A1(n301), .A2(n286), .A3(n117), .A4(n116), .ZN(n300) );
  AOI221_X1 U315 ( .B1(n302), .B2(n289), .C1(n666), .C2(n557), .A(n631), .ZN(
        n301) );
  OAI22_X1 U316 ( .A1(n564), .A2(n161), .B1(n655), .B2(n303), .ZN(n302) );
  NAND4_X1 U317 ( .A1(n196), .A2(n285), .A3(n117), .A4(n116), .ZN(n284) );
  OAI22_X1 U318 ( .A1(n286), .A2(n557), .B1(n287), .B2(n659), .ZN(n285) );
  AOI22_X1 U319 ( .A1(n288), .A2(n289), .B1(n666), .B2(n562), .ZN(n287) );
  OAI221_X1 U320 ( .B1(n607), .B2(n546), .C1(n677), .C2(n550), .A(n387), .ZN(
        N1167) );
  NOR2_X1 U321 ( .A1(n548), .A2(n557), .ZN(n389) );
  AOI221_X1 U322 ( .B1(n652), .B2(n560), .C1(n391), .C2(n392), .A(n393), .ZN(
        n388) );
  OAI221_X1 U323 ( .B1(n622), .B2(n544), .C1(n623), .C2(n550), .A(n227), .ZN(
        N1180) );
  AOI21_X1 U324 ( .B1(n229), .B2(n230), .A(n631), .ZN(n228) );
  OAI221_X1 U325 ( .B1(n593), .B2(n544), .C1(n599), .C2(n550), .A(n414), .ZN(
        N1163) );
  INV_X1 U326 ( .A(n416), .ZN(n635) );
  AOI22_X1 U327 ( .A1(n643), .A2(n557), .B1(n126), .B2(n127), .ZN(n125) );
  AOI21_X1 U328 ( .B1(n573), .B2(n466), .A(n129), .ZN(n126) );
  OAI221_X1 U329 ( .B1(n614), .B2(n543), .C1(n675), .C2(n550), .A(n353), .ZN(
        N1170) );
  OAI22_X1 U330 ( .A1(n355), .A2(n557), .B1(n653), .B2(n356), .ZN(n354) );
  AOI22_X1 U331 ( .A1(n357), .A2(n358), .B1(n507), .B2(n562), .ZN(n356) );
  OAI221_X1 U332 ( .B1(n591), .B2(n543), .C1(n595), .C2(n550), .A(n420), .ZN(
        N1162) );
  OAI211_X1 U333 ( .C1(n553), .C2(n417), .A(n633), .B(n421), .ZN(n420) );
  INV_X1 U334 ( .A(n87), .ZN(n647) );
  INV_X1 U335 ( .A(n89), .ZN(n630) );
  OAI221_X1 U336 ( .B1(n599), .B2(n546), .C1(n603), .C2(n550), .A(n409), .ZN(
        N1164) );
  OAI21_X1 U337 ( .B1(n410), .B2(n411), .A(n633), .ZN(n409) );
  OAI221_X1 U338 ( .B1(n366), .B2(n574), .C1(n530), .C2(n585), .A(n412), .ZN(
        n411) );
  OAI221_X1 U339 ( .B1(n620), .B2(n546), .C1(n621), .C2(n550), .A(n255), .ZN(
        N1178) );
  OAI21_X1 U340 ( .B1(n256), .B2(n257), .A(n196), .ZN(n255) );
  OAI221_X1 U341 ( .B1(n560), .B2(n117), .C1(n116), .C2(n557), .A(n258), .ZN(
        n257) );
  OAI221_X1 U342 ( .B1(n259), .B2(n160), .C1(n161), .C2(n585), .A(n260), .ZN(
        n256) );
  OAI22_X1 U343 ( .A1(n161), .A2(n568), .B1(n655), .B2(n290), .ZN(n288) );
  NAND4_X1 U344 ( .A1(n293), .A2(n294), .A3(n295), .A4(n296), .ZN(n292) );
  NOR3_X1 U345 ( .A1(n273), .A2(n663), .A3(n655), .ZN(n272) );
  OAI21_X1 U346 ( .B1(n586), .B2(n100), .A(n274), .ZN(n273) );
  NAND4_X1 U347 ( .A1(n275), .A2(n276), .A3(n277), .A4(n278), .ZN(n274) );
  OAI211_X1 U348 ( .C1(n624), .C2(n550), .A(n212), .B(n213), .ZN(N1181) );
  AOI22_X1 U350 ( .A1(n551), .A2(n665), .B1(n646), .B2(r1[25]), .ZN(n212) );
  AOI221_X1 U351 ( .B1(n657), .B2(n563), .C1(n565), .C2(n664), .A(n214), .ZN(
        n213) );
  AOI21_X1 U352 ( .B1(n215), .B2(n216), .A(n631), .ZN(n214) );
  OAI211_X1 U353 ( .C1(n625), .C2(n550), .A(n194), .B(n195), .ZN(N1182) );
  AOI22_X1 U354 ( .A1(n551), .A2(n660), .B1(n646), .B2(r1[26]), .ZN(n194) );
  AOI221_X1 U355 ( .B1(n196), .B2(n197), .C1(n573), .C2(n664), .A(n198), .ZN(
        n195) );
  OAI22_X1 U356 ( .A1(n560), .A2(n119), .B1(n199), .B2(n569), .ZN(n198) );
  AOI221_X1 U357 ( .B1(n138), .B2(n654), .C1(n606), .C2(n655), .A(n139), .ZN(
        n137) );
  OAI22_X1 U358 ( .A1(n611), .A2(n100), .B1(n677), .B2(n101), .ZN(n139) );
  NAND2_X1 U359 ( .A1(r2[3]), .A2(n436), .ZN(n85) );
  OAI22_X1 U360 ( .A1(n622), .A2(n529), .B1(n534), .B2(n621), .ZN(n144) );
  AOI22_X1 U361 ( .A1(n604), .A2(n663), .B1(r1[11]), .B2(n656), .ZN(n186) );
  AOI22_X1 U362 ( .A1(n606), .A2(n663), .B1(n656), .B2(n542), .ZN(n162) );
  OAI22_X1 U363 ( .A1(n626), .A2(n550), .B1(n177), .B2(n89), .ZN(N1183) );
  AOI211_X1 U364 ( .C1(n646), .C2(r1[27]), .A(n179), .B(n178), .ZN(n177) );
  OAI22_X1 U365 ( .A1(n472), .A2(n557), .B1(n560), .B2(n118), .ZN(n179) );
  OAI221_X1 U366 ( .B1(n180), .B2(n153), .C1(n154), .C2(n585), .A(n181), .ZN(
        n178) );
  OAI22_X1 U368 ( .A1(n627), .A2(n550), .B1(n148), .B2(n89), .ZN(N1184) );
  NOR2_X1 U369 ( .A1(n149), .A2(n150), .ZN(n148) );
  OAI221_X1 U370 ( .B1(n560), .B2(n472), .C1(n626), .C2(n544), .A(n151), .ZN(
        n150) );
  OAI221_X1 U371 ( .B1(n152), .B2(n153), .C1(n154), .C2(n587), .A(n155), .ZN(
        n149) );
  AOI22_X1 U372 ( .A1(n542), .A2(n652), .B1(n609), .B2(n645), .ZN(n266) );
  AND3_X1 U373 ( .A1(n671), .A2(n670), .A3(r2[3]), .ZN(n440) );
  AOI221_X1 U374 ( .B1(n654), .B2(n217), .C1(n592), .C2(n655), .A(n218), .ZN(
        n216) );
  OAI22_X1 U375 ( .A1(n100), .A2(n603), .B1(n101), .B2(n599), .ZN(n218) );
  NAND4_X1 U376 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(n217) );
  AOI222_X1 U377 ( .A1(n644), .A2(r1[18]), .B1(n604), .B2(n667), .C1(n650), 
        .C2(r1[17]), .ZN(n219) );
  NAND2_X1 U378 ( .A1(n659), .A2(r2[3]), .ZN(n134) );
  NOR2_X1 U379 ( .A1(n182), .A2(n183), .ZN(n180) );
  OAI221_X1 U380 ( .B1(n117), .B2(n591), .C1(n116), .C2(n589), .A(n184), .ZN(
        n183) );
  OAI221_X1 U381 ( .B1(n185), .B2(n160), .C1(n161), .C2(n603), .A(n186), .ZN(
        n182) );
  AOI22_X1 U382 ( .A1(n596), .A2(n666), .B1(n592), .B2(n659), .ZN(n184) );
  INV_X1 U383 ( .A(r1[22]), .ZN(n620) );
  NOR2_X1 U384 ( .A1(n156), .A2(n157), .ZN(n152) );
  OAI221_X1 U385 ( .B1(n117), .B2(n594), .C1(n116), .C2(n591), .A(n158), .ZN(
        n157) );
  OAI221_X1 U386 ( .B1(n159), .B2(n160), .C1(n161), .C2(n605), .A(n162), .ZN(
        n156) );
  AOI22_X1 U387 ( .A1(n601), .A2(n666), .B1(n597), .B2(n659), .ZN(n158) );
  CLKBUF_X1 U388 ( .A(r1[9]), .Z(n601) );
  AOI22_X1 U389 ( .A1(n601), .A2(n663), .B1(n604), .B2(n656), .ZN(n200) );
  AOI22_X1 U390 ( .A1(n654), .A2(n204), .B1(n598), .B2(n655), .ZN(n201) );
  BUF_X1 U391 ( .A(n558), .Z(n562) );
  CLKBUF_X1 U392 ( .A(r1[9]), .Z(n600) );
  INV_X1 U393 ( .A(r1[18]), .ZN(n616) );
  BUF_X1 U394 ( .A(r1[13]), .Z(n608) );
  BUF_X1 U395 ( .A(n559), .Z(n564) );
  BUF_X1 U396 ( .A(n559), .Z(n563) );
  CLKBUF_X1 U397 ( .A(r1[8]), .Z(n597) );
  BUF_X1 U398 ( .A(r1[13]), .Z(n609) );
  CLKBUF_X1 U399 ( .A(r1[8]), .Z(n598) );
  BUF_X1 U400 ( .A(r1[21]), .Z(n617) );
  CLKBUF_X1 U401 ( .A(r1[8]), .Z(n596) );
  BUF_X1 U402 ( .A(n558), .Z(n561) );
  BUF_X1 U403 ( .A(r1[14]), .Z(n612) );
  BUF_X1 U404 ( .A(r1[14]), .Z(n613) );
  INV_X1 U405 ( .A(r2[4]), .ZN(n668) );
  CLKBUF_X1 U406 ( .A(r1[9]), .Z(n602) );
  BUF_X1 U407 ( .A(r1[13]), .Z(n610) );
  BUF_X1 U408 ( .A(r1[21]), .Z(n618) );
  CLKBUF_X1 U409 ( .A(r1[4]), .Z(n583) );
  CLKBUF_X1 U410 ( .A(r1[4]), .Z(n584) );
  OAI221_X1 U411 ( .B1(n547), .B2(n677), .C1(n539), .C2(n607), .A(n252), .ZN(
        n250) );
  AOI22_X1 U412 ( .A1(n604), .A2(n507), .B1(n602), .B2(n653), .ZN(n252) );
  OAI221_X1 U413 ( .B1(n549), .B2(n588), .C1(n539), .C2(n585), .A(n341), .ZN(
        n339) );
  AOI22_X1 U414 ( .A1(n573), .A2(n507), .B1(n565), .B2(n653), .ZN(n341) );
  OAI221_X1 U415 ( .B1(n547), .B2(n591), .C1(n539), .C2(n588), .A(n331), .ZN(
        n329) );
  AOI22_X1 U416 ( .A1(n580), .A2(n507), .B1(n573), .B2(n653), .ZN(n331) );
  OAI221_X1 U417 ( .B1(n548), .B2(n595), .C1(n539), .C2(n591), .A(n321), .ZN(
        n319) );
  AOI22_X1 U418 ( .A1(n586), .A2(n507), .B1(n581), .B2(n653), .ZN(n321) );
  AOI221_X1 U419 ( .B1(n641), .B2(r1[25]), .C1(n457), .C2(r1[26]), .A(n145), 
        .ZN(n142) );
  OAI221_X1 U420 ( .B1(n366), .B2(n599), .C1(n531), .C2(n603), .A(n376), .ZN(
        n375) );
  AOI22_X1 U421 ( .A1(n646), .A2(n600), .B1(n523), .B2(n604), .ZN(n404) );
  NOR2_X1 U422 ( .A1(n405), .A2(n406), .ZN(n402) );
  OAI221_X1 U423 ( .B1(n366), .B2(n585), .C1(n531), .C2(n588), .A(n407), .ZN(
        n406) );
  OAI22_X1 U424 ( .A1(n529), .A2(n675), .B1(n535), .B2(n614), .ZN(n297) );
  OAI22_X1 U425 ( .A1(n529), .A2(n676), .B1(n534), .B2(n673), .ZN(n223) );
  INV_X1 U426 ( .A(r1[15]), .ZN(n675) );
  INV_X1 U427 ( .A(r1[19]), .ZN(n673) );
  AOI221_X1 U428 ( .B1(r1[16]), .B2(n640), .C1(n609), .C2(n650), .A(n280), 
        .ZN(n277) );
  OAI22_X1 U429 ( .A1(n534), .A2(n675), .B1(n532), .B2(n616), .ZN(n280) );
  OAI221_X1 U430 ( .B1(n313), .B2(n270), .C1(n314), .C2(n315), .A(n316), .ZN(
        N1174) );
  AOI22_X1 U431 ( .A1(n646), .A2(r1[18]), .B1(n523), .B2(r1[19]), .ZN(n316) );
  AOI222_X1 U432 ( .A1(n565), .A2(n656), .B1(n552), .B2(n655), .C1(n663), .C2(
        n563), .ZN(n313) );
  NOR4_X1 U433 ( .A1(n317), .A2(n318), .A3(n319), .A4(n320), .ZN(n314) );
  AOI22_X1 U434 ( .A1(r1[18]), .A2(n652), .B1(r1[19]), .B2(n645), .ZN(n173) );
  OAI221_X1 U435 ( .B1(n540), .B2(n676), .C1(n538), .C2(n619), .A(n267), .ZN(
        n261) );
  AOI22_X1 U436 ( .A1(r1[16]), .A2(n639), .B1(r1[17]), .B2(n640), .ZN(n267) );
  INV_X1 U437 ( .A(r1[20]), .ZN(n676) );
  AOI221_X1 U438 ( .B1(r1[16]), .B2(n507), .C1(r1[15]), .C2(n653), .A(n146), 
        .ZN(n141) );
  INV_X1 U439 ( .A(r1[16]), .ZN(n674) );
  OAI221_X1 U440 ( .B1(n335), .B2(n315), .C1(n100), .C2(n557), .A(n336), .ZN(
        N1172) );
  AOI22_X1 U441 ( .A1(n646), .A2(r1[16]), .B1(n523), .B2(r1[17]), .ZN(n336) );
  NOR4_X1 U442 ( .A1(n337), .A2(n338), .A3(n339), .A4(n340), .ZN(n335) );
  OAI221_X1 U443 ( .B1(n241), .B2(n631), .C1(n154), .C2(n557), .A(n242), .ZN(
        N1179) );
  AOI22_X1 U444 ( .A1(n646), .A2(r1[23]), .B1(n523), .B2(r1[24]), .ZN(n242) );
  NOR2_X1 U445 ( .A1(n243), .A2(n244), .ZN(n241) );
  OAI221_X1 U446 ( .B1(n117), .B2(n567), .C1(n560), .C2(n116), .A(n245), .ZN(
        n244) );
  INV_X1 U447 ( .A(r1[11]), .ZN(n607) );
  OAI22_X1 U448 ( .A1(n528), .A2(n619), .B1(n535), .B2(n676), .ZN(n209) );
  AOI22_X1 U449 ( .A1(r1[15]), .A2(n507), .B1(n612), .B2(n653), .ZN(n170) );
  AOI221_X1 U450 ( .B1(r1[17]), .B2(n507), .C1(r1[16]), .C2(n653), .A(n112), 
        .ZN(n103) );
  NAND4_X1 U451 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n204) );
  AOI222_X1 U452 ( .A1(n644), .A2(r1[19]), .B1(n606), .B2(n667), .C1(n650), 
        .C2(r1[18]), .ZN(n205) );
  AOI221_X1 U453 ( .B1(n608), .B2(n507), .C1(n542), .C2(n653), .A(n211), .ZN(
        n206) );
  OAI22_X1 U454 ( .A1(n100), .A2(n599), .B1(n101), .B2(n595), .ZN(n232) );
  NAND4_X1 U455 ( .A1(n233), .A2(n234), .A3(n235), .A4(n236), .ZN(n231) );
  AOI222_X1 U456 ( .A1(n644), .A2(r1[17]), .B1(n601), .B2(n667), .C1(n650), 
        .C2(r1[16]), .ZN(n233) );
  AOI221_X1 U457 ( .B1(r1[20]), .B2(n638), .C1(r1[17]), .C2(n641), .A(n279), 
        .ZN(n278) );
  OAI21_X1 U458 ( .B1(n540), .B2(n673), .A(n100), .ZN(n279) );
  INV_X1 U459 ( .A(r1[27]), .ZN(n625) );
  INV_X1 U460 ( .A(r1[28]), .ZN(n626) );
  CLKBUF_X1 U461 ( .A(r1[1]), .Z(n558) );
  CLKBUF_X1 U462 ( .A(r1[1]), .Z(n559) );
  CLKBUF_X1 U463 ( .A(r1[12]), .Z(n542) );
  BUF_X1 U464 ( .A(n113), .Z(n539) );
  INV_X1 U465 ( .A(n113), .ZN(n648) );
  NAND2_X1 U466 ( .A1(n435), .A2(n433), .ZN(n111) );
  BUF_X1 U467 ( .A(n169), .Z(n524) );
  CLKBUF_X1 U468 ( .A(n169), .Z(n525) );
  CLKBUF_X1 U469 ( .A(n169), .Z(n526) );
  NAND2_X1 U470 ( .A1(n440), .A2(n502), .ZN(n169) );
  OR3_X1 U471 ( .A1(r2[15]), .A2(r2[14]), .A3(r2[13]), .ZN(n451) );
  OAI22_X1 U472 ( .A1(n107), .A2(n623), .B1(n108), .B2(n622), .ZN(n106) );
  INV_X1 U473 ( .A(n494), .ZN(n638) );
  OAI221_X1 U474 ( .B1(n377), .B2(n677), .C1(n167), .C2(n587), .A(n378), .ZN(
        n374) );
  OAI221_X1 U475 ( .B1(n377), .B2(n599), .C1(n560), .C2(n167), .A(n408), .ZN(
        n405) );
  OAI221_X1 U479 ( .B1(n377), .B2(n595), .C1(n167), .C2(n557), .A(n413), .ZN(
        n410) );
  NAND4_X1 U481 ( .A1(n128), .A2(n471), .A3(n443), .A4(n417), .ZN(n377) );
  OAI221_X1 U482 ( .B1(n398), .B2(n399), .C1(n564), .C2(n110), .A(n547), .ZN(
        n396) );
  OAI21_X1 U484 ( .B1(n565), .B2(n110), .A(n549), .ZN(n393) );
  OAI222_X1 U485 ( .A1(n565), .A2(n111), .B1(n383), .B2(n384), .C1(n573), .C2(
        n110), .ZN(n382) );
  OAI222_X1 U486 ( .A1(n579), .A2(n111), .B1(n361), .B2(n362), .C1(n586), .C2(
        n110), .ZN(n360) );
  OAI22_X1 U487 ( .A1(n548), .A2(n605), .B1(n110), .B2(n677), .ZN(n281) );
  OAI22_X1 U489 ( .A1(n110), .A2(n615), .B1(n111), .B2(n674), .ZN(n210) );
  OAI22_X1 U490 ( .A1(n110), .A2(n674), .B1(n111), .B2(n675), .ZN(n224) );
  OAI22_X1 U491 ( .A1(n110), .A2(n675), .B1(n111), .B2(n614), .ZN(n238) );
  OAI22_X1 U492 ( .A1(n110), .A2(n607), .B1(n111), .B2(n605), .ZN(n298) );
  OAI22_X1 U493 ( .A1(n676), .A2(n110), .B1(n111), .B2(n673), .ZN(n145) );
  OAI22_X1 U494 ( .A1(n110), .A2(n619), .B1(n111), .B2(n676), .ZN(n109) );
  NAND2_X1 U495 ( .A1(n642), .A2(r2[3]), .ZN(n527) );
  BUF_X1 U496 ( .A(n114), .Z(n549) );
  BUF_X1 U497 ( .A(n114), .Z(n548) );
  INV_X1 U498 ( .A(n114), .ZN(n636) );
  CLKBUF_X1 U499 ( .A(n124), .Z(n530) );
  AOI221_X1 U500 ( .B1(r1[23]), .B2(n637), .C1(n638), .C2(r1[24]), .A(n223), 
        .ZN(n222) );
  AOI221_X1 U501 ( .B1(r1[18]), .B2(n637), .C1(r1[19]), .C2(n638), .A(n297), 
        .ZN(n296) );
  CLKBUF_X1 U502 ( .A(n171), .Z(n537) );
  CLKBUF_X1 U503 ( .A(n171), .Z(n536) );
  NAND2_X1 U504 ( .A1(n433), .A2(n438), .ZN(n121) );
  NAND2_X1 U505 ( .A1(n436), .A2(n433), .ZN(n417) );
  OAI211_X1 U506 ( .C1(n363), .C2(n677), .A(n513), .B(n365), .ZN(n362) );
  OAI21_X1 U507 ( .B1(n374), .B2(n375), .A(n364), .ZN(n373) );
  OAI211_X1 U508 ( .C1(n363), .C2(n605), .A(n513), .B(n385), .ZN(n384) );
  OAI21_X1 U509 ( .B1(n363), .B2(n603), .A(n513), .ZN(n395) );
  OAI211_X1 U510 ( .C1(n363), .C2(n599), .A(n513), .B(n400), .ZN(n399) );
  OAI211_X1 U511 ( .C1(n552), .C2(n525), .A(n633), .B(n415), .ZN(n414) );
  AOI21_X1 U512 ( .B1(n635), .B2(n526), .A(n650), .ZN(n415) );
  NAND4_X1 U513 ( .A1(n633), .A2(n417), .A3(n167), .A4(n525), .ZN(n426) );
  OAI222_X1 U514 ( .A1(n167), .A2(n603), .B1(n455), .B2(n570), .C1(n526), .C2(
        n605), .ZN(n330) );
  OAI222_X1 U515 ( .A1(n167), .A2(n605), .B1(n455), .B2(n578), .C1(n526), .C2(
        n607), .ZN(n320) );
  OAI222_X1 U516 ( .A1(n167), .A2(n599), .B1(n455), .B2(n560), .C1(n526), .C2(
        n603), .ZN(n340) );
  OAI222_X1 U517 ( .A1(n167), .A2(n595), .B1(n455), .B2(n557), .C1(n526), .C2(
        n599), .ZN(n348) );
  OAI222_X1 U518 ( .A1(n167), .A2(n577), .B1(n377), .B2(n605), .C1(n525), .C2(
        n585), .ZN(n394) );
  OAI222_X1 U519 ( .A1(n167), .A2(n614), .B1(n455), .B2(n595), .C1(n675), .C2(
        n525), .ZN(n264) );
  OAI211_X1 U520 ( .C1(n525), .C2(n677), .A(n291), .B(n309), .ZN(n308) );
  AOI22_X1 U521 ( .A1(n648), .A2(n566), .B1(n359), .B2(n360), .ZN(n357) );
  NOR2_X1 U522 ( .A1(n636), .A2(n648), .ZN(n359) );
  NAND4_X1 U523 ( .A1(n143), .A2(n141), .A3(n142), .A4(n140), .ZN(n138) );
  OAI211_X1 U524 ( .C1(n131), .C2(n132), .A(n630), .B(n647), .ZN(n130) );
  NAND2_X1 U525 ( .A1(n550), .A2(n469), .ZN(n89) );
  NAND2_X1 U526 ( .A1(n643), .A2(n473), .ZN(n107) );
  OAI222_X1 U527 ( .A1(n94), .A2(n557), .B1(n133), .B2(n486), .C1(n560), .C2(
        n134), .ZN(n131) );
  INV_X1 U528 ( .A(n174), .ZN(n637) );
  AOI21_X1 U529 ( .B1(n642), .B2(n560), .A(n129), .ZN(n427) );
  AOI222_X1 U530 ( .A1(n466), .A2(n560), .B1(n128), .B2(n567), .C1(n642), .C2(
        n557), .ZN(n430) );
  AOI22_X1 U531 ( .A1(n580), .A2(n456), .B1(r1[2]), .B2(n642), .ZN(n127) );
  AOI22_X1 U532 ( .A1(n590), .A2(n642), .B1(n592), .B2(n466), .ZN(n407) );
  AOI22_X1 U533 ( .A1(n586), .A2(n642), .B1(r1[6]), .B2(n466), .ZN(n412) );
  AOI22_X1 U534 ( .A1(n573), .A2(n642), .B1(n586), .B2(n128), .ZN(n424) );
  AOI222_X1 U535 ( .A1(n585), .A2(n642), .B1(n591), .B2(n128), .C1(n589), .C2(
        n466), .ZN(n419) );
  AOI22_X1 U536 ( .A1(n604), .A2(n642), .B1(n606), .B2(n466), .ZN(n376) );
  NOR2_X1 U537 ( .A1(n466), .A2(n642), .ZN(n128) );
  NAND2_X1 U538 ( .A1(n642), .A2(r2[3]), .ZN(n114) );
  CLKBUF_X1 U539 ( .A(n124), .Z(n531) );
  NAND2_X1 U540 ( .A1(n442), .A2(n433), .ZN(n124) );
  NAND2_X1 U541 ( .A1(n634), .A2(n351), .ZN(n403) );
  NAND2_X1 U542 ( .A1(n351), .A2(n642), .ZN(n172) );
  BUF_X2 U543 ( .A(n108), .Z(n534) );
  NAND2_X1 U544 ( .A1(n500), .A2(n651), .ZN(n108) );
  OR4_X2 U545 ( .A1(r2[27]), .A2(r2[26]), .A3(r2[29]), .A4(r2[28]), .ZN(n449)
         );
  NAND2_X1 U546 ( .A1(n515), .A2(n351), .ZN(n175) );
  AOI211_X1 U547 ( .C1(n422), .C2(n417), .A(n644), .B(n650), .ZN(n421) );
  AOI22_X1 U548 ( .A1(n565), .A2(n644), .B1(n573), .B2(n651), .ZN(n408) );
  AOI22_X1 U549 ( .A1(n644), .A2(n561), .B1(r1[2]), .B2(n651), .ZN(n413) );
  AOI222_X1 U550 ( .A1(n579), .A2(n651), .B1(n602), .B2(n515), .C1(n571), .C2(
        n644), .ZN(n401) );
  AOI221_X1 U551 ( .B1(n612), .B2(n644), .C1(n606), .C2(n652), .A(n281), .ZN(
        n276) );
  AOI222_X1 U552 ( .A1(n590), .A2(n651), .B1(n606), .B2(n515), .C1(r1[5]), 
        .C2(n644), .ZN(n386) );
  AOI222_X1 U553 ( .A1(n596), .A2(n651), .B1(n609), .B2(n515), .C1(r1[7]), 
        .C2(n644), .ZN(n368) );
  AOI22_X1 U554 ( .A1(n590), .A2(n644), .B1(n592), .B2(n651), .ZN(n378) );
  AOI222_X1 U555 ( .A1(n608), .A2(n644), .B1(n586), .B2(n667), .C1(n542), .C2(
        n650), .ZN(n293) );
  AOI222_X1 U556 ( .A1(n644), .A2(r1[22]), .B1(n612), .B2(n667), .C1(n650), 
        .C2(n617), .ZN(n140) );
  AOI222_X1 U557 ( .A1(r1[23]), .A2(n644), .B1(r1[15]), .B2(n667), .C1(r1[22]), 
        .C2(n650), .ZN(n102) );
  NAND2_X1 U558 ( .A1(n514), .A2(r2[3]), .ZN(n113) );
  NAND2_X1 U559 ( .A1(n466), .A2(n351), .ZN(n174) );
  CLKBUF_X1 U560 ( .A(n390), .Z(n541) );
  OAI22_X1 U561 ( .A1(n92), .A2(n486), .B1(n94), .B2(n560), .ZN(n91) );
  AOI211_X1 U562 ( .C1(n565), .C2(n465), .A(n90), .B(n91), .ZN(n88) );
  INV_X1 U563 ( .A(r2[0]), .ZN(n672) );
  AOI22_X1 U564 ( .A1(n427), .A2(n428), .B1(n553), .B2(n649), .ZN(n425) );
  OAI211_X1 U565 ( .C1(n564), .C2(n530), .A(n632), .B(n125), .ZN(n123) );
  OAI221_X1 U566 ( .B1(n536), .B2(n611), .C1(n532), .C2(n614), .A(n332), .ZN(
        n328) );
  OAI221_X1 U567 ( .B1(n537), .B2(n614), .C1(n533), .C2(n675), .A(n322), .ZN(
        n318) );
  OAI221_X1 U568 ( .B1(n536), .B2(n677), .C1(n532), .C2(n611), .A(n342), .ZN(
        n338) );
  OAI221_X1 U569 ( .B1(n537), .B2(n607), .C1(n533), .C2(n677), .A(n350), .ZN(
        n346) );
  OAI221_X1 U570 ( .B1(n561), .B2(n366), .C1(n565), .C2(n531), .A(n423), .ZN(
        n422) );
  AOI22_X1 U571 ( .A1(n565), .A2(n650), .B1(r1[6]), .B2(n649), .ZN(n400) );
  OAI221_X1 U572 ( .B1(n536), .B2(n673), .C1(n532), .C2(n676), .A(n253), .ZN(
        n249) );
  OAI222_X1 U573 ( .A1(n366), .A2(n565), .B1(n530), .B2(n573), .C1(n129), .C2(
        n419), .ZN(n418) );
  OAI221_X1 U574 ( .B1(n537), .B2(n616), .C1(n533), .C2(n673), .A(n266), .ZN(
        n262) );
  AOI22_X1 U575 ( .A1(n580), .A2(n650), .B1(n597), .B2(n649), .ZN(n385) );
  OAI221_X1 U576 ( .B1(n622), .B2(n536), .C1(n623), .C2(n532), .A(n173), .ZN(
        n164) );
  AOI211_X1 U577 ( .C1(n97), .C2(n96), .A(n657), .B(n664), .ZN(n95) );
  OAI221_X1 U578 ( .B1(n537), .B2(n675), .C1(n533), .C2(n674), .A(n311), .ZN(
        n306) );
  AOI22_X1 U579 ( .A1(n590), .A2(n650), .B1(n604), .B2(n649), .ZN(n365) );
  OAI221_X1 U580 ( .B1(n536), .B2(n621), .C1(n622), .C2(n533), .A(n192), .ZN(
        n188) );
  INV_X1 U581 ( .A(n171), .ZN(n641) );
  NAND2_X1 U582 ( .A1(n473), .A2(n649), .ZN(n171) );
  OAI211_X1 U583 ( .C1(n552), .C2(n111), .A(n541), .B(n485), .ZN(n397) );
  OAI211_X1 U584 ( .C1(n388), .C2(n389), .A(n541), .B(n485), .ZN(n387) );
  OAI22_X1 U585 ( .A1(n283), .A2(n599), .B1(n539), .B2(n603), .ZN(n282) );
  OAI22_X1 U586 ( .A1(n539), .A2(n614), .B1(n547), .B2(n675), .ZN(n211) );
  OAI22_X1 U587 ( .A1(n539), .A2(n611), .B1(n547), .B2(n614), .ZN(n225) );
  OAI22_X1 U588 ( .A1(n539), .A2(n677), .B1(n549), .B2(n611), .ZN(n239) );
  OAI22_X1 U589 ( .A1(n539), .A2(n599), .B1(n114), .B2(n603), .ZN(n299) );
  OAI22_X1 U590 ( .A1(n539), .A2(n615), .B1(n114), .B2(n616), .ZN(n146) );
  OAI22_X1 U591 ( .A1(n539), .A2(n616), .B1(n114), .B2(n673), .ZN(n112) );
  INV_X1 U592 ( .A(n523), .ZN(n550) );
  INV_X1 U593 ( .A(r1[2]), .ZN(n566) );
  INV_X1 U594 ( .A(r1[2]), .ZN(n567) );
  INV_X1 U595 ( .A(r1[2]), .ZN(n568) );
  INV_X1 U596 ( .A(r1[2]), .ZN(n569) );
  INV_X1 U597 ( .A(r1[2]), .ZN(n570) );
  CLKBUF_X1 U598 ( .A(r1[3]), .Z(n571) );
  CLKBUF_X1 U599 ( .A(r1[3]), .Z(n572) );
  INV_X1 U600 ( .A(n571), .ZN(n574) );
  INV_X1 U601 ( .A(n571), .ZN(n575) );
  INV_X1 U602 ( .A(n571), .ZN(n576) );
  INV_X1 U603 ( .A(n572), .ZN(n577) );
  INV_X1 U604 ( .A(r1[3]), .ZN(n578) );
  INV_X1 U605 ( .A(r1[5]), .ZN(n587) );
  INV_X1 U606 ( .A(r1[5]), .ZN(n588) );
  INV_X1 U607 ( .A(r1[5]), .ZN(n589) );
  INV_X1 U608 ( .A(r1[6]), .ZN(n591) );
  INV_X1 U609 ( .A(r1[7]), .ZN(n593) );
  INV_X1 U610 ( .A(r1[7]), .ZN(n594) );
  INV_X1 U611 ( .A(r1[7]), .ZN(n595) );
  INV_X1 U612 ( .A(r1[10]), .ZN(n605) );
  INV_X1 U613 ( .A(r1[17]), .ZN(n615) );
  INV_X1 U614 ( .A(n618), .ZN(n619) );
  INV_X1 U615 ( .A(r1[23]), .ZN(n621) );
  INV_X1 U616 ( .A(r1[24]), .ZN(n622) );
  INV_X1 U617 ( .A(r1[25]), .ZN(n623) );
  INV_X1 U618 ( .A(r1[26]), .ZN(n624) );
  INV_X1 U619 ( .A(r1[29]), .ZN(n627) );
  INV_X1 U620 ( .A(r1[30]), .ZN(n628) );
  INV_X2 U621 ( .A(n524), .ZN(n644) );
  INV_X2 U622 ( .A(n417), .ZN(n651) );
  INV_X2 U623 ( .A(n168), .ZN(n667) );
endmodule


module shifter_dx_nbit32 ( r1, r2, log, data_out );
  input [31:0] r1;
  input [31:0] r2;
  output [31:0] data_out;
  input log;
  wire   N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069,
         N2070, N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079,
         N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089,
         N2090, N2091, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803;

  DLH_X1 \data_out_reg[31]  ( .G(1'b1), .D(N2091), .Q(data_out[31]) );
  DLH_X1 \data_out_reg[30]  ( .G(1'b1), .D(N2090), .Q(data_out[30]) );
  DLH_X1 \data_out_reg[29]  ( .G(1'b1), .D(N2089), .Q(data_out[29]) );
  DLH_X1 \data_out_reg[28]  ( .G(1'b1), .D(N2088), .Q(data_out[28]) );
  DLH_X1 \data_out_reg[27]  ( .G(1'b1), .D(N2087), .Q(data_out[27]) );
  DLH_X1 \data_out_reg[26]  ( .G(1'b1), .D(N2086), .Q(data_out[26]) );
  DLH_X1 \data_out_reg[25]  ( .G(1'b1), .D(N2085), .Q(data_out[25]) );
  DLH_X1 \data_out_reg[24]  ( .G(1'b1), .D(N2084), .Q(data_out[24]) );
  DLH_X1 \data_out_reg[23]  ( .G(1'b1), .D(N2083), .Q(data_out[23]) );
  DLH_X1 \data_out_reg[22]  ( .G(1'b1), .D(N2082), .Q(data_out[22]) );
  DLH_X1 \data_out_reg[21]  ( .G(1'b1), .D(N2081), .Q(data_out[21]) );
  DLH_X1 \data_out_reg[20]  ( .G(1'b1), .D(N2080), .Q(data_out[20]) );
  DLH_X1 \data_out_reg[19]  ( .G(1'b1), .D(N2079), .Q(data_out[19]) );
  DLH_X1 \data_out_reg[18]  ( .G(1'b1), .D(N2078), .Q(data_out[18]) );
  DLH_X1 \data_out_reg[17]  ( .G(1'b1), .D(N2077), .Q(data_out[17]) );
  DLH_X1 \data_out_reg[16]  ( .G(1'b1), .D(N2076), .Q(data_out[16]) );
  DLH_X1 \data_out_reg[15]  ( .G(1'b1), .D(N2075), .Q(data_out[15]) );
  DLH_X1 \data_out_reg[14]  ( .G(1'b1), .D(N2074), .Q(data_out[14]) );
  DLH_X1 \data_out_reg[13]  ( .G(1'b1), .D(N2073), .Q(data_out[13]) );
  DLH_X1 \data_out_reg[12]  ( .G(1'b1), .D(N2072), .Q(data_out[12]) );
  DLH_X1 \data_out_reg[11]  ( .G(1'b1), .D(N2071), .Q(data_out[11]) );
  DLH_X1 \data_out_reg[10]  ( .G(1'b1), .D(N2070), .Q(data_out[10]) );
  DLH_X1 \data_out_reg[9]  ( .G(1'b1), .D(N2069), .Q(data_out[9]) );
  DLH_X1 \data_out_reg[8]  ( .G(1'b1), .D(N2068), .Q(data_out[8]) );
  DLH_X1 \data_out_reg[7]  ( .G(1'b1), .D(N2067), .Q(data_out[7]) );
  DLH_X1 \data_out_reg[6]  ( .G(1'b1), .D(N2066), .Q(data_out[6]) );
  DLH_X1 \data_out_reg[5]  ( .G(1'b1), .D(N2065), .Q(data_out[5]) );
  DLH_X1 \data_out_reg[4]  ( .G(1'b1), .D(N2064), .Q(data_out[4]) );
  DLH_X1 \data_out_reg[3]  ( .G(1'b1), .D(N2063), .Q(data_out[3]) );
  DLH_X1 \data_out_reg[2]  ( .G(1'b1), .D(N2062), .Q(data_out[2]) );
  DLH_X1 \data_out_reg[1]  ( .G(1'b1), .D(N2061), .Q(data_out[1]) );
  DLH_X1 \data_out_reg[0]  ( .G(1'b1), .D(N2060), .Q(data_out[0]) );
  NAND2_X2 U367 ( .A1(n481), .A2(n489), .ZN(n284) );
  NAND2_X2 U392 ( .A1(n482), .A2(n652), .ZN(n196) );
  AND3_X2 U408 ( .A1(n774), .A2(n798), .A3(r2[4]), .ZN(n479) );
  NAND3_X1 U524 ( .A1(n123), .A2(n124), .A3(n125), .ZN(n121) );
  NAND3_X1 U525 ( .A1(n746), .A2(n135), .A3(n626), .ZN(n131) );
  NAND3_X1 U526 ( .A1(n659), .A2(n661), .A3(n140), .ZN(n139) );
  NAND3_X1 U527 ( .A1(n656), .A2(n662), .A3(r1[25]), .ZN(n156) );
  NAND3_X1 U528 ( .A1(n179), .A2(n180), .A3(n181), .ZN(N2080) );
  NAND3_X1 U529 ( .A1(n761), .A2(n185), .A3(n186), .ZN(n184) );
  NAND3_X1 U530 ( .A1(n187), .A2(n188), .A3(n189), .ZN(n182) );
  NAND3_X1 U531 ( .A1(n203), .A2(n204), .A3(n205), .ZN(n199) );
  NAND3_X1 U533 ( .A1(n314), .A2(n315), .A3(n316), .ZN(N2070) );
  NAND3_X1 U534 ( .A1(n373), .A2(n374), .A3(n375), .ZN(n369) );
  NAND3_X1 U535 ( .A1(n419), .A2(n420), .A3(n421), .ZN(N2063) );
  NAND3_X1 U536 ( .A1(n425), .A2(n427), .A3(n426), .ZN(n424) );
  NAND3_X1 U537 ( .A1(n435), .A2(n436), .A3(n437), .ZN(N2062) );
  NAND3_X1 U538 ( .A1(n763), .A2(n105), .A3(log), .ZN(n158) );
  NAND3_X1 U539 ( .A1(n450), .A2(n751), .A3(n451), .ZN(N2061) );
  NAND3_X1 U540 ( .A1(n372), .A2(n387), .A3(n371), .ZN(n334) );
  INV_X1 U3 ( .A(n780), .ZN(n553) );
  INV_X2 U4 ( .A(n227), .ZN(n781) );
  AND3_X2 U5 ( .A1(r2[0]), .A2(n774), .A3(r2[4]), .ZN(n481) );
  OAI222_X1 U6 ( .A1(n695), .A2(n646), .B1(n697), .B2(n644), .C1(n656), .C2(
        n801), .ZN(n292) );
  OAI221_X1 U7 ( .B1(n654), .B2(n665), .C1(n196), .C2(n676), .A(n467), .ZN(
        n463) );
  OAI222_X1 U8 ( .A1(n646), .A2(n691), .B1(n695), .B2(n644), .C1(n655), .C2(
        n679), .ZN(n310) );
  NOR3_X1 U9 ( .A1(n796), .A2(r2[1]), .A3(n795), .ZN(n482) );
  BUF_X1 U10 ( .A(n498), .Z(n652) );
  NOR3_X1 U11 ( .A1(r2[1]), .A2(r2[2]), .A3(n795), .ZN(n483) );
  BUF_X1 U12 ( .A(n608), .Z(n653) );
  INV_X1 U13 ( .A(n624), .ZN(n230) );
  NAND2_X1 U14 ( .A1(n482), .A2(n606), .ZN(n227) );
  OAI222_X1 U15 ( .A1(n699), .A2(n285), .B1(n412), .B2(n605), .C1(n697), .C2(
        n284), .ZN(n410) );
  OR2_X1 U16 ( .A1(n297), .A2(n775), .ZN(n620) );
  AND2_X1 U17 ( .A1(n575), .A2(n576), .ZN(n174) );
  INV_X1 U18 ( .A(n566), .ZN(n106) );
  OR2_X2 U19 ( .A1(n582), .A2(n334), .ZN(n566) );
  INV_X1 U20 ( .A(n571), .ZN(n98) );
  BUF_X1 U21 ( .A(n176), .Z(n607) );
  AND3_X1 U22 ( .A1(n397), .A2(n396), .A3(n395), .ZN(n554) );
  OR3_X1 U23 ( .A1(n361), .A2(n363), .A3(n362), .ZN(n555) );
  OR3_X1 U24 ( .A1(n310), .A2(n312), .A3(n311), .ZN(n556) );
  OR3_X1 U25 ( .A1(n465), .A2(n464), .A3(n466), .ZN(n557) );
  OR3_X1 U26 ( .A1(n292), .A2(n293), .A3(n294), .ZN(n558) );
  OR3_X1 U27 ( .A1(n415), .A2(n416), .A3(n414), .ZN(n559) );
  AND2_X1 U28 ( .A1(n304), .A2(n301), .ZN(n560) );
  OR3_X1 U29 ( .A1(r2[17]), .A2(r2[18]), .A3(r2[16]), .ZN(n561) );
  OR3_X1 U30 ( .A1(r2[24]), .A2(r2[25]), .A3(r2[23]), .ZN(n562) );
  OR2_X1 U31 ( .A1(n798), .A2(r2[4]), .ZN(n563) );
  AND2_X1 U32 ( .A1(n594), .A2(n593), .ZN(n564) );
  OR2_X1 U33 ( .A1(n753), .A2(n756), .ZN(n565) );
  NOR2_X1 U34 ( .A1(n281), .A2(n565), .ZN(n280) );
  BUF_X2 U35 ( .A(n168), .Z(n646) );
  BUF_X2 U36 ( .A(n197), .Z(n644) );
  AOI221_X1 U37 ( .B1(r1[20]), .B2(n788), .C1(r1[19]), .C2(n107), .A(n791), 
        .ZN(n236) );
  NOR2_X1 U38 ( .A1(n413), .A2(n559), .ZN(n412) );
  NOR3_X1 U39 ( .A1(n567), .A2(n568), .A3(n569), .ZN(n441) );
  NAND3_X1 U40 ( .A1(n622), .A2(n621), .A3(n623), .ZN(n567) );
  AND2_X1 U41 ( .A1(n760), .A2(n683), .ZN(n568) );
  AND2_X1 U42 ( .A1(n790), .A2(n680), .ZN(n569) );
  CLKBUF_X1 U43 ( .A(n763), .Z(n570) );
  NAND2_X1 U44 ( .A1(n479), .A2(n489), .ZN(n270) );
  NAND2_X1 U45 ( .A1(n479), .A2(n497), .ZN(n285) );
  NAND2_X2 U46 ( .A1(n479), .A2(n491), .ZN(n249) );
  AND2_X1 U47 ( .A1(n491), .A2(n653), .ZN(n571) );
  BUF_X1 U48 ( .A(n490), .Z(n606) );
  AND3_X2 U49 ( .A1(n477), .A2(n476), .A3(n407), .ZN(n371) );
  NAND3_X1 U50 ( .A1(n207), .A2(n215), .A3(n107), .ZN(n572) );
  NAND3_X1 U51 ( .A1(n207), .A2(n215), .A3(n107), .ZN(n573) );
  INV_X1 U52 ( .A(n145), .ZN(n574) );
  AND2_X1 U53 ( .A1(n499), .A2(n652), .ZN(n625) );
  BUF_X1 U54 ( .A(n490), .Z(n650) );
  NOR2_X1 U55 ( .A1(n647), .A2(n563), .ZN(n490) );
  NAND2_X1 U56 ( .A1(n185), .A2(n186), .ZN(n575) );
  INV_X1 U57 ( .A(n157), .ZN(n576) );
  INV_X1 U58 ( .A(n582), .ZN(n185) );
  NAND2_X1 U59 ( .A1(n398), .A2(n554), .ZN(n394) );
  AOI221_X1 U60 ( .B1(n688), .B2(n788), .C1(r1[20]), .C2(n107), .A(n791), .ZN(
        n221) );
  NAND2_X1 U61 ( .A1(n306), .A2(n560), .ZN(n299) );
  OR2_X1 U62 ( .A1(n98), .A2(n673), .ZN(n577) );
  OR2_X1 U63 ( .A1(n101), .A2(n803), .ZN(n578) );
  NAND3_X1 U64 ( .A1(n577), .A2(n578), .A3(n298), .ZN(N2071) );
  BUF_X1 U65 ( .A(n127), .Z(n579) );
  AND2_X1 U66 ( .A1(n715), .A2(n600), .ZN(n580) );
  AND2_X1 U67 ( .A1(n725), .A2(n601), .ZN(n581) );
  NOR3_X1 U68 ( .A1(n580), .A2(n581), .A3(n749), .ZN(n110) );
  NAND2_X1 U69 ( .A1(n278), .A2(n564), .ZN(N2072) );
  OR3_X2 U70 ( .A1(n755), .A2(n767), .A3(n296), .ZN(n582) );
  AOI21_X2 U71 ( .B1(n582), .B2(n736), .A(n264), .ZN(n163) );
  AND2_X1 U72 ( .A1(n680), .A2(n600), .ZN(n583) );
  AND2_X1 U73 ( .A1(n624), .A2(n776), .ZN(n584) );
  NOR3_X1 U74 ( .A1(n225), .A2(n584), .A3(n583), .ZN(n224) );
  CLKBUF_X3 U75 ( .A(n572), .Z(n654) );
  BUF_X1 U76 ( .A(n145), .Z(n649) );
  OAI221_X1 U77 ( .B1(n654), .B2(n668), .C1(n196), .C2(n800), .A(n417), .ZN(
        n413) );
  NAND2_X1 U78 ( .A1(n369), .A2(n268), .ZN(n585) );
  NAND2_X1 U79 ( .A1(n737), .A2(n370), .ZN(n586) );
  AND3_X1 U80 ( .A1(n585), .A2(n586), .A3(n751), .ZN(n368) );
  NAND2_X1 U81 ( .A1(n770), .A2(n700), .ZN(n587) );
  NAND2_X1 U82 ( .A1(n214), .A2(n377), .ZN(n588) );
  NAND2_X1 U83 ( .A1(n759), .A2(n704), .ZN(n589) );
  AND3_X1 U84 ( .A1(n587), .A2(n588), .A3(n589), .ZN(n374) );
  BUF_X2 U85 ( .A(n490), .Z(n651) );
  NOR2_X1 U86 ( .A1(n463), .A2(n557), .ZN(n462) );
  OR2_X1 U87 ( .A1(n691), .A2(n285), .ZN(n590) );
  OR2_X1 U88 ( .A1(n462), .A2(n605), .ZN(n591) );
  OR2_X1 U89 ( .A1(n802), .A2(n284), .ZN(n592) );
  NAND3_X1 U90 ( .A1(n590), .A2(n591), .A3(n592), .ZN(n460) );
  OR2_X1 U91 ( .A1(n98), .A2(n803), .ZN(n593) );
  OR2_X1 U92 ( .A1(n101), .A2(n676), .ZN(n594) );
  INV_X1 U93 ( .A(n601), .ZN(n101) );
  NOR2_X1 U94 ( .A1(n360), .A2(n555), .ZN(n359) );
  AND2_X1 U95 ( .A1(n790), .A2(n694), .ZN(n595) );
  AND2_X1 U96 ( .A1(n760), .A2(n696), .ZN(n596) );
  NOR3_X1 U97 ( .A1(n595), .A2(n596), .A3(n358), .ZN(n357) );
  OAI222_X1 U98 ( .A1(n802), .A2(n285), .B1(n487), .B2(n605), .C1(n799), .C2(
        n284), .ZN(n485) );
  OAI221_X1 U99 ( .B1(n654), .B2(n664), .C1(n196), .C2(n803), .A(n496), .ZN(
        n492) );
  NOR2_X1 U100 ( .A1(n309), .A2(n556), .ZN(n308) );
  OR2_X1 U101 ( .A1(n707), .A2(n247), .ZN(n597) );
  OR2_X1 U102 ( .A1(n308), .A2(n222), .ZN(n598) );
  OR2_X1 U103 ( .A1(n712), .A2(n249), .ZN(n599) );
  NAND3_X1 U104 ( .A1(n597), .A2(n598), .A3(n599), .ZN(n305) );
  NAND2_X1 U105 ( .A1(n249), .A2(n247), .ZN(n222) );
  AND2_X1 U106 ( .A1(n284), .A2(n285), .ZN(n488) );
  INV_X1 U107 ( .A(n284), .ZN(n770) );
  INV_X1 U108 ( .A(n285), .ZN(n759) );
  BUF_X1 U109 ( .A(n641), .Z(n642) );
  INV_X2 U110 ( .A(n98), .ZN(n600) );
  AND2_X4 U111 ( .A1(n651), .A2(n491), .ZN(n601) );
  OR4_X2 U112 ( .A1(r2[7]), .A2(r2[6]), .A3(r2[8]), .A4(r2[9]), .ZN(n505) );
  OR4_X1 U113 ( .A1(r2[27]), .A2(r2[26]), .A3(r2[29]), .A4(r2[28]), .ZN(n506)
         );
  NOR2_X1 U114 ( .A1(n507), .A2(n561), .ZN(n502) );
  NOR2_X1 U115 ( .A1(n291), .A2(n558), .ZN(n290) );
  OR2_X1 U116 ( .A1(n712), .A2(n247), .ZN(n602) );
  OR2_X1 U117 ( .A1(n290), .A2(n222), .ZN(n603) );
  OR2_X1 U118 ( .A1(n718), .A2(n249), .ZN(n604) );
  NAND3_X1 U119 ( .A1(n602), .A2(n603), .A3(n604), .ZN(n288) );
  OR4_X1 U120 ( .A1(r2[20]), .A2(r2[19]), .A3(r2[22]), .A4(r2[21]), .ZN(n507)
         );
  NAND2_X2 U121 ( .A1(n480), .A2(n651), .ZN(n247) );
  INV_X1 U122 ( .A(n625), .ZN(n145) );
  OR2_X2 U123 ( .A1(n222), .A2(n582), .ZN(n605) );
  NOR3_X1 U124 ( .A1(r2[0]), .A2(r2[4]), .A3(n647), .ZN(n608) );
  NOR3_X1 U125 ( .A1(r2[0]), .A2(r2[4]), .A3(n647), .ZN(n498) );
  INV_X2 U126 ( .A(n793), .ZN(n640) );
  INV_X1 U127 ( .A(n227), .ZN(n609) );
  NAND2_X1 U128 ( .A1(n608), .A2(n483), .ZN(n177) );
  OR2_X1 U129 ( .A1(n713), .A2(n285), .ZN(n610) );
  OR2_X1 U130 ( .A1(n359), .A2(n605), .ZN(n611) );
  OR2_X1 U131 ( .A1(n706), .A2(n284), .ZN(n612) );
  NAND3_X1 U132 ( .A1(n610), .A2(n611), .A3(n612), .ZN(n358) );
  OAI221_X1 U133 ( .B1(n654), .B2(n671), .C1(n196), .C2(n799), .A(n364), .ZN(
        n360) );
  OR2_X1 U134 ( .A1(n98), .A2(n667), .ZN(n613) );
  OR2_X1 U135 ( .A1(n101), .A2(n668), .ZN(n614) );
  NAND3_X1 U136 ( .A1(n613), .A2(n614), .A3(n383), .ZN(N2065) );
  NAND2_X1 U137 ( .A1(n123), .A2(n384), .ZN(n615) );
  NAND2_X1 U138 ( .A1(n385), .A2(n776), .ZN(n616) );
  AND3_X1 U139 ( .A1(n615), .A2(n616), .A3(n751), .ZN(n383) );
  NOR3_X1 U140 ( .A1(n601), .A2(n571), .A3(n648), .ZN(n123) );
  AND2_X1 U141 ( .A1(r1[9]), .A2(n600), .ZN(n617) );
  AND2_X1 U142 ( .A1(n333), .A2(n745), .ZN(n618) );
  AND2_X1 U143 ( .A1(n758), .A2(n776), .ZN(n619) );
  NOR3_X1 U144 ( .A1(n617), .A2(n618), .A3(n619), .ZN(n328) );
  NAND2_X1 U145 ( .A1(n105), .A2(n752), .ZN(n297) );
  OR2_X1 U146 ( .A1(n695), .A2(n285), .ZN(n621) );
  OR2_X1 U147 ( .A1(n443), .A2(n605), .ZN(n622) );
  OR2_X1 U148 ( .A1(n691), .A2(n284), .ZN(n623) );
  OAI221_X1 U149 ( .B1(n654), .B2(n666), .C1(n196), .C2(n679), .A(n448), .ZN(
        n444) );
  AND2_X4 U150 ( .A1(n480), .A2(n653), .ZN(n624) );
  BUF_X1 U151 ( .A(n99), .Z(n648) );
  BUF_X1 U152 ( .A(n153), .Z(n641) );
  AND3_X1 U153 ( .A1(n643), .A2(n645), .A3(n196), .ZN(n207) );
  INV_X1 U154 ( .A(n643), .ZN(n779) );
  INV_X1 U155 ( .A(n645), .ZN(n791) );
  NOR3_X1 U156 ( .A1(r2[1]), .A2(r2[3]), .A3(n796), .ZN(n497) );
  NOR3_X1 U157 ( .A1(r2[2]), .A2(r2[3]), .A3(n797), .ZN(n489) );
  NOR3_X1 U158 ( .A1(r2[2]), .A2(r2[3]), .A3(r2[1]), .ZN(n491) );
  NOR3_X1 U159 ( .A1(n796), .A2(r2[3]), .A3(n797), .ZN(n499) );
  NAND2_X1 U160 ( .A1(n650), .A2(n483), .ZN(n176) );
  NOR3_X1 U161 ( .A1(n786), .A2(n574), .A3(n150), .ZN(n626) );
  OR2_X1 U162 ( .A1(n733), .A2(n372), .ZN(n627) );
  OR2_X1 U163 ( .A1(n722), .A2(n387), .ZN(n628) );
  NAND3_X1 U164 ( .A1(n627), .A2(n628), .A3(n388), .ZN(n384) );
  NAND2_X1 U165 ( .A1(r1[7]), .A2(n600), .ZN(n629) );
  NAND2_X1 U166 ( .A1(n762), .A2(n736), .ZN(n630) );
  INV_X1 U167 ( .A(n355), .ZN(n631) );
  AND3_X1 U168 ( .A1(n629), .A2(n630), .A3(n631), .ZN(n354) );
  OR2_X1 U169 ( .A1(n802), .A2(n247), .ZN(n632) );
  OR2_X1 U170 ( .A1(n691), .A2(n249), .ZN(n633) );
  NAND3_X1 U171 ( .A1(n632), .A2(n633), .A3(n393), .ZN(n389) );
  NAND2_X1 U172 ( .A1(r1[7]), .A2(n778), .ZN(n634) );
  NAND2_X1 U173 ( .A1(n680), .A2(n792), .ZN(n635) );
  INV_X1 U174 ( .A(n399), .ZN(n636) );
  AND3_X1 U175 ( .A1(n634), .A2(n635), .A3(n636), .ZN(n398) );
  INV_X1 U176 ( .A(n196), .ZN(n792) );
  NOR2_X1 U177 ( .A1(n506), .A2(n562), .ZN(n503) );
  NAND2_X1 U178 ( .A1(n770), .A2(n698), .ZN(n637) );
  NAND2_X1 U179 ( .A1(n214), .A2(n394), .ZN(n638) );
  NAND2_X1 U180 ( .A1(n759), .A2(n700), .ZN(n639) );
  AND3_X1 U181 ( .A1(n637), .A2(n638), .A3(n639), .ZN(n393) );
  NOR2_X1 U182 ( .A1(n105), .A2(n100), .ZN(n162) );
  INV_X1 U183 ( .A(r1[24]), .ZN(n699) );
  INV_X1 U184 ( .A(n119), .ZN(n761) );
  INV_X1 U185 ( .A(n215), .ZN(n780) );
  NOR2_X1 U186 ( .A1(n781), .A2(n624), .ZN(n215) );
  NAND2_X1 U187 ( .A1(n202), .A2(n207), .ZN(n119) );
  INV_X1 U188 ( .A(n116), .ZN(n742) );
  INV_X1 U189 ( .A(n282), .ZN(n756) );
  NOR3_X1 U190 ( .A1(n769), .A2(n768), .A3(n758), .ZN(n282) );
  NOR2_X1 U191 ( .A1(n222), .A2(n582), .ZN(n214) );
  NOR2_X1 U192 ( .A1(n620), .A2(n566), .ZN(n157) );
  OAI21_X1 U193 ( .B1(n163), .B2(n620), .A(n751), .ZN(n116) );
  INV_X1 U194 ( .A(n318), .ZN(n776) );
  INV_X1 U195 ( .A(n607), .ZN(n787) );
  NOR2_X1 U196 ( .A1(n780), .A2(n222), .ZN(n202) );
  OAI21_X1 U197 ( .B1(n620), .B2(n404), .A(n751), .ZN(n423) );
  INV_X1 U198 ( .A(n247), .ZN(n790) );
  INV_X1 U199 ( .A(n334), .ZN(n763) );
  INV_X1 U200 ( .A(n123), .ZN(n775) );
  INV_X1 U201 ( .A(n343), .ZN(n748) );
  INV_X1 U202 ( .A(n268), .ZN(n747) );
  INV_X1 U203 ( .A(n454), .ZN(n766) );
  INV_X1 U204 ( .A(n730), .ZN(n733) );
  INV_X1 U205 ( .A(n138), .ZN(n794) );
  INV_X1 U206 ( .A(n137), .ZN(n789) );
  INV_X1 U207 ( .A(n108), .ZN(n788) );
  AOI211_X1 U208 ( .C1(n761), .C2(n199), .A(n201), .B(n183), .ZN(n200) );
  OAI22_X1 U209 ( .A1(n722), .A2(n646), .B1(n733), .B2(n644), .ZN(n201) );
  INV_X1 U210 ( .A(n319), .ZN(n769) );
  NAND2_X1 U211 ( .A1(n123), .A2(n736), .ZN(n318) );
  INV_X1 U212 ( .A(n332), .ZN(n768) );
  AOI21_X1 U213 ( .B1(n222), .B2(n112), .A(n116), .ZN(n223) );
  AOI21_X1 U214 ( .B1(n150), .B2(n112), .A(n749), .ZN(n141) );
  NAND4_X1 U215 ( .A1(n319), .A2(n332), .A3(n366), .A4(n488), .ZN(n296) );
  AOI21_X1 U216 ( .B1(n296), .B2(n736), .A(n264), .ZN(n271) );
  INV_X1 U217 ( .A(n366), .ZN(n758) );
  AOI22_X1 U218 ( .A1(n730), .A2(n770), .B1(n737), .B2(n759), .ZN(n301) );
  OAI21_X1 U219 ( .B1(n764), .B2(n772), .A(n737), .ZN(n404) );
  NAND2_X1 U220 ( .A1(n123), .A2(n105), .ZN(n454) );
  AOI21_X1 U221 ( .B1(n134), .B2(n264), .A(n162), .ZN(n343) );
  NAND2_X1 U222 ( .A1(n134), .A2(n570), .ZN(n244) );
  AOI22_X1 U223 ( .A1(n794), .A2(n736), .B1(n117), .B2(n118), .ZN(n114) );
  OAI22_X1 U224 ( .A1(n733), .A2(n657), .B1(n784), .B2(n722), .ZN(n117) );
  INV_X1 U225 ( .A(n249), .ZN(n760) );
  INV_X1 U226 ( .A(n387), .ZN(n762) );
  NAND2_X1 U227 ( .A1(n753), .A2(n244), .ZN(n268) );
  NOR3_X1 U228 ( .A1(n773), .A2(n764), .A3(n765), .ZN(n477) );
  INV_X1 U229 ( .A(n162), .ZN(n751) );
  INV_X1 U230 ( .A(n161), .ZN(n749) );
  AOI21_X1 U231 ( .B1(n127), .B2(n134), .A(n162), .ZN(n161) );
  INV_X1 U232 ( .A(n408), .ZN(n773) );
  INV_X1 U233 ( .A(n372), .ZN(n771) );
  INV_X1 U234 ( .A(n476), .ZN(n772) );
  CLKBUF_X1 U235 ( .A(n108), .Z(n655) );
  CLKBUF_X1 U236 ( .A(n137), .Z(n658) );
  CLKBUF_X1 U237 ( .A(n138), .Z(n661) );
  CLKBUF_X1 U238 ( .A(n108), .Z(n656) );
  CLKBUF_X1 U239 ( .A(n137), .Z(n659) );
  CLKBUF_X1 U240 ( .A(n138), .Z(n662) );
  CLKBUF_X1 U241 ( .A(n108), .Z(n657) );
  CLKBUF_X1 U242 ( .A(n138), .Z(n663) );
  CLKBUF_X1 U243 ( .A(n137), .Z(n660) );
  INV_X1 U244 ( .A(n174), .ZN(n745) );
  INV_X1 U245 ( .A(n386), .ZN(n765) );
  NAND2_X1 U246 ( .A1(n229), .A2(n230), .ZN(n228) );
  INV_X1 U247 ( .A(n455), .ZN(n764) );
  INV_X1 U248 ( .A(n144), .ZN(n746) );
  INV_X1 U249 ( .A(n118), .ZN(n743) );
  INV_X1 U250 ( .A(n648), .ZN(n774) );
  NOR3_X1 U251 ( .A1(n797), .A2(n796), .A3(n795), .ZN(n480) );
  NOR2_X1 U252 ( .A1(n297), .A2(n775), .ZN(n134) );
  INV_X1 U253 ( .A(n726), .ZN(n722) );
  NOR2_X1 U254 ( .A1(n576), .A2(n740), .ZN(n112) );
  NOR3_X1 U255 ( .A1(n797), .A2(r2[2]), .A3(n795), .ZN(n478) );
  INV_X1 U256 ( .A(n703), .ZN(n700) );
  AOI222_X1 U257 ( .A1(n768), .A2(n710), .B1(n758), .B2(n704), .C1(n769), .C2(
        n700), .ZN(n418) );
  AOI222_X1 U258 ( .A1(n787), .A2(n700), .B1(n779), .B2(n710), .C1(n791), .C2(
        n704), .ZN(n240) );
  INV_X1 U259 ( .A(n690), .ZN(n691) );
  AOI222_X1 U260 ( .A1(n624), .A2(n729), .B1(n792), .B2(n715), .C1(n609), .C2(
        n724), .ZN(n239) );
  INV_X1 U261 ( .A(n693), .ZN(n695) );
  NOR2_X1 U262 ( .A1(n738), .A2(n763), .ZN(n264) );
  OAI221_X1 U263 ( .B1(n685), .B2(n270), .C1(n682), .C2(n287), .A(n500), .ZN(
        n484) );
  AOI222_X1 U264 ( .A1(n768), .A2(n696), .B1(n758), .B2(n692), .C1(n769), .C2(
        n687), .ZN(n500) );
  AOI211_X1 U265 ( .C1(n783), .C2(n129), .A(n566), .B(n119), .ZN(n126) );
  INV_X1 U266 ( .A(n124), .ZN(n783) );
  OAI21_X1 U267 ( .B1(n119), .B2(n576), .A(n184), .ZN(n118) );
  INV_X1 U268 ( .A(n675), .ZN(n676) );
  INV_X1 U269 ( .A(n678), .ZN(n679) );
  AOI22_X1 U270 ( .A1(n761), .A2(n157), .B1(n123), .B2(n125), .ZN(n144) );
  OAI221_X1 U271 ( .B1(n283), .B2(n770), .C1(n737), .C2(n284), .A(n285), .ZN(
        n281) );
  AOI22_X1 U272 ( .A1(n286), .A2(n270), .B1(n755), .B2(n733), .ZN(n283) );
  OAI22_X1 U273 ( .A1(n726), .A2(n287), .B1(n288), .B2(n767), .ZN(n286) );
  NOR3_X1 U274 ( .A1(n332), .A2(n738), .A3(n244), .ZN(n331) );
  AOI211_X1 U275 ( .C1(n106), .C2(n305), .A(n307), .B(n264), .ZN(n306) );
  OAI21_X1 U276 ( .B1(n761), .B2(n738), .A(n163), .ZN(n127) );
  NAND2_X1 U277 ( .A1(n480), .A2(n481), .ZN(n105) );
  AOI22_X1 U278 ( .A1(n733), .A2(n779), .B1(n644), .B2(n198), .ZN(n195) );
  OAI22_X1 U279 ( .A1(n199), .A2(n791), .B1(n646), .B2(n724), .ZN(n198) );
  AOI22_X1 U280 ( .A1(r1[28]), .A2(n767), .B1(n726), .B2(n755), .ZN(n304) );
  NAND2_X1 U281 ( .A1(n479), .A2(n499), .ZN(n366) );
  NAND2_X1 U282 ( .A1(n482), .A2(n479), .ZN(n407) );
  NAND2_X1 U283 ( .A1(n478), .A2(n479), .ZN(n386) );
  INV_X1 U284 ( .A(r2[1]), .ZN(n797) );
  INV_X1 U285 ( .A(r2[2]), .ZN(n796) );
  INV_X1 U286 ( .A(n684), .ZN(n685) );
  AOI22_X1 U287 ( .A1(n771), .A2(n700), .B1(n762), .B2(n698), .ZN(n473) );
  AOI22_X1 U288 ( .A1(n288), .A2(n106), .B1(n755), .B2(n728), .ZN(n289) );
  AOI22_X1 U289 ( .A1(n789), .A2(n710), .B1(r1[26]), .B2(n794), .ZN(n166) );
  AOI22_X1 U290 ( .A1(n771), .A2(n704), .B1(n762), .B2(n700), .ZN(n456) );
  AOI22_X1 U291 ( .A1(n793), .A2(n710), .B1(n787), .B2(n715), .ZN(n204) );
  AOI221_X1 U292 ( .B1(n696), .B2(n794), .C1(n694), .C2(n788), .A(n206), .ZN(
        n205) );
  OAI211_X1 U293 ( .C1(n740), .C2(n646), .A(n169), .B(n170), .ZN(N2081) );
  AOI22_X1 U294 ( .A1(n171), .A2(n761), .B1(n112), .B2(n119), .ZN(n169) );
  AOI21_X1 U295 ( .B1(n172), .B2(n173), .A(n174), .ZN(n171) );
  INV_X1 U296 ( .A(n741), .ZN(n736) );
  OAI211_X1 U297 ( .C1(n101), .C2(n703), .A(n141), .B(n142), .ZN(N2084) );
  OAI211_X1 U298 ( .C1(n733), .C2(n145), .A(n146), .B(n147), .ZN(n143) );
  AOI222_X1 U299 ( .A1(n789), .A2(n725), .B1(r1[27]), .B2(n788), .C1(n794), 
        .C2(n715), .ZN(n147) );
  OAI211_X1 U300 ( .C1(n101), .C2(n679), .A(n265), .B(n266), .ZN(N2073) );
  AOI211_X1 U301 ( .C1(n267), .C2(n268), .A(n269), .B(n162), .ZN(n266) );
  OAI22_X1 U302 ( .A1(n739), .A2(n270), .B1(n271), .B2(n620), .ZN(n269) );
  OAI22_X1 U303 ( .A1(n739), .A2(n98), .B1(n648), .B2(n100), .ZN(N2091) );
  NAND2_X1 U304 ( .A1(n480), .A2(n479), .ZN(n455) );
  NAND2_X1 U305 ( .A1(n481), .A2(n483), .ZN(n372) );
  NOR2_X1 U306 ( .A1(n780), .A2(n211), .ZN(n193) );
  NOR2_X1 U307 ( .A1(n740), .A2(n282), .ZN(n307) );
  OAI21_X1 U308 ( .B1(n605), .B2(n244), .A(n211), .ZN(n229) );
  NAND4_X1 U309 ( .A1(n210), .A2(n214), .A3(n553), .A4(n570), .ZN(n213) );
  AOI21_X1 U310 ( .B1(n737), .B2(n406), .A(n162), .ZN(n405) );
  OAI21_X1 U311 ( .B1(n297), .B2(n407), .A(n408), .ZN(n406) );
  OAI211_X1 U312 ( .C1(n303), .C2(n754), .A(n285), .B(n284), .ZN(n302) );
  INV_X1 U313 ( .A(n304), .ZN(n754) );
  AND3_X1 U314 ( .A1(n305), .A2(n287), .A3(n270), .ZN(n303) );
  NAND2_X1 U315 ( .A1(n479), .A2(n483), .ZN(n387) );
  AOI22_X1 U316 ( .A1(n793), .A2(n715), .B1(n787), .B2(n723), .ZN(n187) );
  AOI221_X1 U317 ( .B1(n700), .B2(n789), .C1(n698), .C2(n794), .A(n190), .ZN(
        n189) );
  OAI211_X1 U318 ( .C1(n113), .C2(n744), .A(n114), .B(n115), .ZN(N2087) );
  INV_X1 U319 ( .A(n112), .ZN(n744) );
  OAI211_X1 U320 ( .C1(n740), .C2(n657), .A(n109), .B(n110), .ZN(N2088) );
  NOR2_X1 U321 ( .A1(n743), .A2(n733), .ZN(n111) );
  NAND4_X1 U322 ( .A1(n131), .A2(n751), .A3(n132), .A4(n133), .ZN(N2085) );
  OAI221_X1 U323 ( .B1(n98), .B2(n733), .C1(n740), .C2(n101), .A(n102), .ZN(
        N2090) );
  BUF_X1 U324 ( .A(n731), .Z(n729) );
  BUF_X1 U325 ( .A(n732), .Z(n728) );
  NAND4_X1 U326 ( .A1(n120), .A2(n121), .A3(n751), .A4(n122), .ZN(N2086) );
  OAI21_X1 U327 ( .B1(n126), .B2(n579), .A(n128), .ZN(n120) );
  BUF_X1 U328 ( .A(n731), .Z(n730) );
  INV_X1 U329 ( .A(n186), .ZN(n753) );
  BUF_X1 U330 ( .A(n732), .Z(n727) );
  INV_X1 U331 ( .A(n391), .ZN(n750) );
  OAI222_X1 U332 ( .A1(n699), .A2(n247), .B1(n335), .B2(n222), .C1(n702), .C2(
        n249), .ZN(n333) );
  NOR4_X1 U333 ( .A1(n336), .A2(n337), .A3(n338), .A4(n339), .ZN(n335) );
  OAI22_X1 U334 ( .A1(n802), .A2(n230), .B1(n799), .B2(n227), .ZN(n382) );
  INV_X1 U335 ( .A(n719), .ZN(n715) );
  NOR4_X1 U336 ( .A1(n492), .A2(n493), .A3(n494), .A4(n495), .ZN(n487) );
  OAI222_X1 U337 ( .A1(n660), .A2(n667), .B1(n649), .B2(n668), .C1(n661), .C2(
        n666), .ZN(n495) );
  OAI222_X1 U338 ( .A1(n658), .A2(n802), .B1(n649), .B2(n691), .C1(n662), .C2(
        n799), .ZN(n253) );
  OAI222_X1 U339 ( .A1(n658), .A2(n803), .B1(n649), .B2(n676), .C1(n662), .C2(
        n673), .ZN(n363) );
  OAI222_X1 U340 ( .A1(n717), .A2(n319), .B1(n722), .B2(n366), .C1(n733), .C2(
        n332), .ZN(n365) );
  OAI222_X1 U341 ( .A1(n711), .A2(n319), .B1(n717), .B2(n366), .C1(n722), .C2(
        n332), .ZN(n376) );
  OAI222_X1 U342 ( .A1(n699), .A2(n319), .B1(n701), .B2(n366), .C1(n706), .C2(
        n332), .ZN(n428) );
  OAI222_X1 U343 ( .A1(n646), .A2(n685), .B1(n644), .B2(n799), .C1(n657), .C2(
        n673), .ZN(n349) );
  OAI222_X1 U344 ( .A1(n318), .A2(n319), .B1(n244), .B2(n757), .C1(n98), .C2(
        n672), .ZN(n317) );
  INV_X1 U345 ( .A(n307), .ZN(n757) );
  OAI222_X1 U346 ( .A1(n658), .A2(n800), .B1(n649), .B2(n682), .C1(n662), .C2(
        n801), .ZN(n312) );
  OAI222_X1 U347 ( .A1(n659), .A2(n679), .B1(n649), .B2(n801), .C1(n663), .C2(
        n676), .ZN(n339) );
  OAI222_X1 U348 ( .A1(n659), .A2(n799), .B1(n649), .B2(n802), .C1(n663), .C2(
        n685), .ZN(n262) );
  NOR4_X1 U349 ( .A1(n444), .A2(n445), .A3(n446), .A4(n447), .ZN(n443) );
  OAI222_X1 U350 ( .A1(n659), .A2(n669), .B1(n649), .B2(n670), .C1(n663), .C2(
        n668), .ZN(n447) );
  OAI222_X1 U351 ( .A1(n722), .A2(n408), .B1(n733), .B2(n407), .C1(n716), .C2(
        n386), .ZN(n438) );
  OAI222_X1 U352 ( .A1(n660), .A2(n668), .B1(n649), .B2(n669), .C1(n661), .C2(
        n667), .ZN(n466) );
  NOR3_X1 U353 ( .A1(n410), .A2(n409), .A3(n411), .ZN(n403) );
  OAI22_X1 U354 ( .A1(n802), .A2(n249), .B1(n799), .B2(n247), .ZN(n411) );
  OAI221_X1 U355 ( .B1(n695), .B2(n270), .C1(n691), .C2(n287), .A(n418), .ZN(
        n409) );
  OAI222_X1 U356 ( .A1(n717), .A2(n285), .B1(n347), .B2(n605), .C1(n712), .C2(
        n284), .ZN(n345) );
  NOR4_X1 U357 ( .A1(n348), .A2(n349), .A3(n350), .A4(n351), .ZN(n347) );
  OAI222_X1 U358 ( .A1(n660), .A2(n676), .B1(n649), .B2(n679), .C1(n661), .C2(
        n803), .ZN(n351) );
  OAI222_X1 U359 ( .A1(n697), .A2(n646), .B1(n699), .B2(n644), .C1(n655), .C2(
        n800), .ZN(n274) );
  OAI222_X1 U360 ( .A1(n646), .A2(n682), .B1(n644), .B2(n685), .C1(n656), .C2(
        n672), .ZN(n361) );
  OAI222_X1 U361 ( .A1(n646), .A2(n799), .B1(n644), .B2(n802), .C1(n655), .C2(
        n803), .ZN(n337) );
  OAI222_X1 U362 ( .A1(n646), .A2(n803), .B1(n644), .B2(n676), .C1(n656), .C2(
        n667), .ZN(n445) );
  OAI222_X1 U363 ( .A1(n646), .A2(n672), .B1(n644), .B2(n673), .C1(n656), .C2(
        n665), .ZN(n493) );
  OAI222_X1 U364 ( .A1(n646), .A2(n673), .B1(n644), .B2(n803), .C1(n655), .C2(
        n666), .ZN(n464) );
  OAI222_X1 U365 ( .A1(n699), .A2(n646), .B1(n701), .B2(n644), .C1(n656), .C2(
        n682), .ZN(n260) );
  OAI222_X1 U366 ( .A1(n646), .A2(n802), .B1(n691), .B2(n644), .C1(n657), .C2(
        n676), .ZN(n323) );
  OAI222_X1 U368 ( .A1(n702), .A2(n646), .B1(n707), .B2(n644), .C1(n657), .C2(
        n685), .ZN(n251) );
  OAI222_X1 U369 ( .A1(n703), .A2(n247), .B1(n321), .B2(n222), .C1(n706), .C2(
        n249), .ZN(n320) );
  NOR4_X1 U370 ( .A1(n322), .A2(n323), .A3(n324), .A4(n325), .ZN(n321) );
  OAI222_X1 U371 ( .A1(n659), .A2(n801), .B1(n649), .B2(n800), .C1(n663), .C2(
        n679), .ZN(n325) );
  OAI222_X1 U372 ( .A1(n722), .A2(n249), .B1(n716), .B2(n247), .C1(n272), .C2(
        n605), .ZN(n267) );
  NOR4_X1 U373 ( .A1(n273), .A2(n274), .A3(n275), .A4(n276), .ZN(n272) );
  OAI222_X1 U374 ( .A1(n660), .A2(n685), .B1(n649), .B2(n799), .C1(n661), .C2(
        n682), .ZN(n276) );
  AOI22_X1 U375 ( .A1(n609), .A2(n692), .B1(n624), .B2(n696), .ZN(n340) );
  AOI22_X1 U376 ( .A1(n609), .A2(n710), .B1(n624), .B2(n715), .ZN(n263) );
  AOI22_X1 U377 ( .A1(n609), .A2(n686), .B1(n624), .B2(n692), .ZN(n352) );
  AOI22_X1 U378 ( .A1(n609), .A2(n704), .B1(n624), .B2(n710), .ZN(n277) );
  AOI22_X1 U379 ( .A1(n609), .A2(n696), .B1(n624), .B2(n698), .ZN(n326) );
  AOI22_X1 U380 ( .A1(n781), .A2(n698), .B1(n624), .B2(n700), .ZN(n313) );
  AOI22_X1 U381 ( .A1(n609), .A2(n715), .B1(n624), .B2(n723), .ZN(n255) );
  OAI222_X1 U382 ( .A1(n660), .A2(n682), .B1(n145), .B2(n685), .C1(n661), .C2(
        n800), .ZN(n294) );
  OAI222_X1 U383 ( .A1(n646), .A2(n679), .B1(n644), .B2(n801), .C1(n657), .C2(
        n669), .ZN(n414) );
  OAI222_X1 U384 ( .A1(n658), .A2(n671), .B1(n649), .B2(n672), .C1(n662), .C2(
        n670), .ZN(n416) );
  AOI221_X1 U385 ( .B1(n704), .B2(n789), .C1(n700), .C2(n794), .A(n178), .ZN(
        n172) );
  OAI22_X1 U386 ( .A1(n714), .A2(n649), .B1(n717), .B2(n642), .ZN(n178) );
  OAI221_X1 U387 ( .B1(n784), .B2(n718), .C1(n722), .C2(n656), .A(n130), .ZN(
        n124) );
  AOI22_X1 U388 ( .A1(n789), .A2(n736), .B1(n794), .B2(n728), .ZN(n130) );
  OAI221_X1 U389 ( .B1(n799), .B2(n270), .C1(n685), .C2(n287), .A(n468), .ZN(
        n459) );
  AOI222_X1 U390 ( .A1(n768), .A2(n698), .B1(n758), .B2(n696), .C1(n769), .C2(
        n693), .ZN(n468) );
  OAI221_X1 U391 ( .B1(n474), .B2(n334), .C1(n718), .C2(n407), .A(n475), .ZN(
        n471) );
  AOI22_X1 U393 ( .A1(n772), .A2(n723), .B1(n773), .B2(n710), .ZN(n475) );
  NOR3_X1 U394 ( .A1(n485), .A2(n484), .A3(n486), .ZN(n474) );
  OAI22_X1 U395 ( .A1(n800), .A2(n249), .B1(n247), .B2(n801), .ZN(n486) );
  OAI221_X1 U396 ( .B1(n697), .B2(n270), .C1(n695), .C2(n287), .A(n392), .ZN(
        n390) );
  AOI222_X1 U397 ( .A1(n768), .A2(r1[28]), .B1(n758), .B2(n710), .C1(n769), 
        .C2(n704), .ZN(n392) );
  OAI221_X1 U398 ( .B1(n457), .B2(n334), .C1(n722), .C2(n407), .A(n458), .ZN(
        n452) );
  AOI22_X1 U399 ( .A1(n772), .A2(n727), .B1(n773), .B2(n715), .ZN(n458) );
  NOR3_X1 U400 ( .A1(n459), .A2(n460), .A3(n461), .ZN(n457) );
  OAI22_X1 U401 ( .A1(n682), .A2(n249), .B1(n247), .B2(n800), .ZN(n461) );
  OAI221_X1 U402 ( .B1(n706), .B2(n270), .C1(n702), .C2(n287), .A(n353), .ZN(
        n344) );
  AOI222_X1 U403 ( .A1(n768), .A2(n736), .B1(n758), .B2(n729), .C1(n769), .C2(
        n724), .ZN(n353) );
  AOI22_X1 U404 ( .A1(n781), .A2(n700), .B1(n624), .B2(n704), .ZN(n295) );
  OAI221_X1 U405 ( .B1(n784), .B2(n699), .C1(n655), .C2(n702), .A(n167), .ZN(
        n164) );
  AOI22_X1 U406 ( .A1(n793), .A2(n727), .B1(n787), .B2(n736), .ZN(n167) );
  NOR3_X1 U407 ( .A1(n119), .A2(n582), .A3(n158), .ZN(n125) );
  OAI21_X1 U409 ( .B1(n371), .B2(n297), .A(n386), .ZN(n385) );
  OAI211_X1 U410 ( .C1(n722), .C2(n287), .A(n271), .B(n289), .ZN(n279) );
  OAI221_X1 U411 ( .B1(n98), .B2(n666), .C1(n101), .C2(n667), .A(n400), .ZN(
        N2064) );
  OAI21_X1 U412 ( .B1(n401), .B2(n402), .A(n123), .ZN(n400) );
  OAI222_X1 U413 ( .A1(n722), .A2(n372), .B1(n733), .B2(n386), .C1(n716), .C2(
        n387), .ZN(n402) );
  OAI221_X1 U414 ( .B1(n750), .B2(n403), .C1(n297), .C2(n404), .A(n405), .ZN(
        n401) );
  AOI221_X1 U415 ( .B1(n134), .B2(n299), .C1(n300), .C2(n282), .A(n162), .ZN(
        n298) );
  AOI21_X1 U416 ( .B1(n301), .B2(n302), .A(n753), .ZN(n300) );
  OAI221_X1 U417 ( .B1(n98), .B2(n799), .C1(n101), .C2(n802), .A(n191), .ZN(
        N2079) );
  AOI221_X1 U418 ( .B1(n128), .B2(n192), .C1(n193), .C2(n777), .A(n162), .ZN(
        n191) );
  INV_X1 U419 ( .A(n194), .ZN(n777) );
  OAI21_X1 U420 ( .B1(n200), .B2(n566), .A(n163), .ZN(n192) );
  OAI221_X1 U421 ( .B1(n98), .B2(n722), .C1(n733), .C2(n101), .A(n103), .ZN(
        N2089) );
  OAI21_X1 U422 ( .B1(n104), .B2(n752), .A(n776), .ZN(n103) );
  OAI221_X1 U423 ( .B1(n733), .B2(n660), .C1(n722), .C2(n661), .A(n139), .ZN(
        n135) );
  OAI22_X1 U424 ( .A1(n788), .A2(n711), .B1(n655), .B2(n716), .ZN(n140) );
  NOR2_X1 U425 ( .A1(n158), .A2(n775), .ZN(n186) );
  OAI22_X1 U426 ( .A1(n658), .A2(n699), .B1(n649), .B2(n701), .ZN(n206) );
  OAI22_X1 U427 ( .A1(n708), .A2(n145), .B1(n714), .B2(n642), .ZN(n190) );
  OAI22_X1 U428 ( .A1(n98), .A2(n665), .B1(n318), .B2(n407), .ZN(n422) );
  OAI221_X1 U429 ( .B1(n743), .B2(n159), .C1(n98), .C2(n695), .A(n160), .ZN(
        N2082) );
  NOR2_X1 U430 ( .A1(n164), .A2(n165), .ZN(n159) );
  AOI21_X1 U431 ( .B1(n696), .B2(n601), .A(n749), .ZN(n160) );
  OAI221_X1 U432 ( .B1(n722), .B2(n642), .C1(n719), .C2(n145), .A(n166), .ZN(
        n165) );
  OAI221_X1 U433 ( .B1(n747), .B2(n341), .C1(n98), .C2(n670), .A(n342), .ZN(
        N2068) );
  AOI21_X1 U434 ( .B1(r1[9]), .B2(n601), .A(n748), .ZN(n342) );
  NOR3_X1 U435 ( .A1(n344), .A2(n345), .A3(n346), .ZN(n341) );
  OAI22_X1 U436 ( .A1(n699), .A2(n249), .B1(n697), .B2(n247), .ZN(n346) );
  AOI22_X1 U437 ( .A1(n779), .A2(n716), .B1(n232), .B2(n644), .ZN(n231) );
  OAI22_X1 U438 ( .A1(r1[27]), .A2(n646), .B1(n233), .B2(n234), .ZN(n232) );
  OAI221_X1 U439 ( .B1(n659), .B2(n695), .C1(n663), .C2(n691), .A(n236), .ZN(
        n233) );
  OAI21_X1 U440 ( .B1(n334), .B2(n297), .A(n158), .ZN(n391) );
  INV_X1 U441 ( .A(n713), .ZN(n710) );
  INV_X1 U442 ( .A(n707), .ZN(n704) );
  OAI22_X1 U443 ( .A1(n722), .A2(n145), .B1(n574), .B2(n154), .ZN(n152) );
  AOI22_X1 U444 ( .A1(n155), .A2(n658), .B1(n789), .B2(n715), .ZN(n154) );
  OAI221_X1 U445 ( .B1(n655), .B2(n708), .C1(n662), .C2(n713), .A(n156), .ZN(
        n155) );
  OAI22_X1 U446 ( .A1(n782), .A2(n779), .B1(n644), .B2(n724), .ZN(n216) );
  INV_X1 U447 ( .A(n217), .ZN(n782) );
  OAI22_X1 U448 ( .A1(r1[28]), .A2(n646), .B1(n218), .B2(n219), .ZN(n217) );
  INV_X1 U449 ( .A(n681), .ZN(n682) );
  INV_X1 U450 ( .A(r2[3]), .ZN(n795) );
  OAI211_X1 U451 ( .C1(n101), .C2(n685), .A(n223), .B(n224), .ZN(N2077) );
  AOI221_X1 U452 ( .B1(n226), .B2(n227), .C1(n609), .C2(n733), .A(n228), .ZN(
        n225) );
  OAI211_X1 U453 ( .C1(n101), .C2(n801), .A(n742), .B(n256), .ZN(N2074) );
  OAI222_X1 U454 ( .A1(n722), .A2(n247), .B1(n258), .B2(n222), .C1(n733), .C2(
        n249), .ZN(n257) );
  NOR4_X1 U455 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(n258) );
  OAI211_X1 U456 ( .C1(n101), .C2(n699), .A(n141), .B(n148), .ZN(N2083) );
  NOR3_X1 U457 ( .A1(n150), .A2(n144), .A3(n151), .ZN(n149) );
  OAI211_X1 U458 ( .C1(n101), .C2(n799), .A(n208), .B(n209), .ZN(N2078) );
  AOI221_X1 U459 ( .B1(n210), .B2(n193), .C1(n609), .C2(n776), .A(n162), .ZN(
        n209) );
  OAI211_X1 U460 ( .C1(n202), .C2(n740), .A(n213), .B(n163), .ZN(n212) );
  NOR4_X1 U461 ( .A1(n505), .A2(r2[30]), .A3(r2[5]), .A4(r2[31]), .ZN(n504) );
  NOR4_X1 U462 ( .A1(n508), .A2(r2[10]), .A3(r2[12]), .A4(r2[11]), .ZN(n501)
         );
  NAND2_X1 U463 ( .A1(n737), .A2(n752), .ZN(n100) );
  AOI22_X1 U464 ( .A1(n790), .A2(n686), .B1(n760), .B2(n692), .ZN(n373) );
  AOI221_X1 U465 ( .B1(n755), .B2(n698), .C1(n767), .C2(n696), .A(n376), .ZN(
        n375) );
  BUF_X1 U466 ( .A(r1[22]), .Z(n692) );
  BUF_X1 U467 ( .A(r1[22]), .Z(n693) );
  BUF_X1 U468 ( .A(n720), .Z(n723) );
  BUF_X1 U469 ( .A(n720), .Z(n724) );
  BUF_X1 U470 ( .A(n721), .Z(n726) );
  BUF_X1 U471 ( .A(r1[18]), .Z(n683) );
  OR3_X1 U472 ( .A1(r2[15]), .A2(r2[14]), .A3(r2[13]), .ZN(n508) );
  BUF_X1 U473 ( .A(n721), .Z(n725) );
  BUF_X1 U474 ( .A(r1[18]), .Z(n684) );
  AOI222_X1 U475 ( .A1(n771), .A2(n715), .B1(n773), .B2(n729), .C1(n765), .C2(
        n725), .ZN(n420) );
  AOI211_X1 U476 ( .C1(r1[4]), .C2(n601), .A(n422), .B(n423), .ZN(n421) );
  AOI22_X1 U477 ( .A1(n762), .A2(n710), .B1(n424), .B2(n268), .ZN(n419) );
  BUF_X1 U478 ( .A(r1[14]), .Z(n677) );
  OR3_X1 U479 ( .A1(n158), .A2(n775), .A3(n605), .ZN(n211) );
  BUF_X1 U480 ( .A(r1[13]), .Z(n674) );
  BUF_X1 U481 ( .A(r1[22]), .Z(n694) );
  BUF_X1 U482 ( .A(r1[14]), .Z(n678) );
  BUF_X1 U483 ( .A(r1[13]), .Z(n675) );
  BUF_X1 U484 ( .A(r1[30]), .Z(n731) );
  BUF_X1 U485 ( .A(r1[30]), .Z(n732) );
  AOI22_X1 U486 ( .A1(n680), .A2(n781), .B1(n624), .B2(n683), .ZN(n417) );
  AOI22_X1 U487 ( .A1(n674), .A2(n781), .B1(n678), .B2(n624), .ZN(n496) );
  INV_X1 U488 ( .A(r1[19]), .ZN(n799) );
  INV_X1 U489 ( .A(r1[20]), .ZN(n802) );
  INV_X1 U490 ( .A(r1[16]), .ZN(n800) );
  AOI221_X1 U491 ( .B1(n778), .B2(n684), .C1(r1[19]), .C2(n788), .A(n243), 
        .ZN(n242) );
  OAI22_X1 U492 ( .A1(n662), .A2(n802), .B1(n658), .B2(n691), .ZN(n243) );
  AOI221_X1 U493 ( .B1(r1[5]), .B2(n778), .C1(r1[15]), .C2(n792), .A(n434), 
        .ZN(n433) );
  OAI22_X1 U494 ( .A1(n230), .A2(n682), .B1(n227), .B2(n800), .ZN(n434) );
  OAI22_X1 U495 ( .A1(n799), .A2(n230), .B1(n227), .B2(n685), .ZN(n399) );
  INV_X1 U496 ( .A(r1[15]), .ZN(n801) );
  INV_X1 U497 ( .A(r1[12]), .ZN(n803) );
  OAI221_X1 U498 ( .B1(n659), .B2(n697), .C1(n663), .C2(n695), .A(n221), .ZN(
        n218) );
  OAI221_X1 U499 ( .B1(n454), .B2(n469), .C1(n318), .C2(n105), .A(n470), .ZN(
        N2060) );
  NOR2_X1 U500 ( .A1(n471), .A2(n472), .ZN(n469) );
  OAI221_X1 U501 ( .B1(n705), .B2(n386), .C1(n733), .C2(n455), .A(n473), .ZN(
        n472) );
  AOI21_X1 U502 ( .B1(n356), .B2(n357), .A(n747), .ZN(n355) );
  AOI221_X1 U503 ( .B1(n755), .B2(n700), .C1(n767), .C2(n698), .A(n365), .ZN(
        n356) );
  OAI211_X1 U504 ( .C1(n101), .C2(n669), .A(n367), .B(n368), .ZN(N2066) );
  OAI21_X1 U505 ( .B1(n371), .B2(n620), .A(n372), .ZN(n370) );
  OAI211_X1 U506 ( .C1(n101), .C2(n800), .A(n742), .B(n245), .ZN(N2075) );
  OAI222_X1 U507 ( .A1(n733), .A2(n247), .B1(n248), .B2(n222), .C1(n738), .C2(
        n249), .ZN(n246) );
  NOR4_X1 U508 ( .A1(n250), .A2(n251), .A3(n252), .A4(n253), .ZN(n248) );
  OAI211_X1 U509 ( .C1(n101), .C2(n682), .A(n223), .B(n237), .ZN(N2076) );
  NAND4_X1 U510 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(n238) );
  NAND4_X1 U511 ( .A1(n378), .A2(n379), .A3(n380), .A4(n381), .ZN(n377) );
  AOI222_X1 U512 ( .A1(r1[10]), .A2(n794), .B1(r1[12]), .B2(n574), .C1(r1[11]), 
        .C2(n789), .ZN(n378) );
  AOI222_X1 U513 ( .A1(r1[9]), .A2(n788), .B1(n681), .B2(n779), .C1(r1[16]), 
        .C2(n791), .ZN(n380) );
  NAND4_X1 U514 ( .A1(n430), .A2(n431), .A3(n432), .A4(n433), .ZN(n429) );
  AOI222_X1 U515 ( .A1(r1[7]), .A2(n794), .B1(r1[9]), .B2(n574), .C1(r1[8]), 
        .C2(n789), .ZN(n430) );
  AOI222_X1 U516 ( .A1(r1[6]), .A2(n788), .B1(n677), .B2(n779), .C1(n675), 
        .C2(n791), .ZN(n432) );
  AOI222_X1 U517 ( .A1(r1[9]), .A2(n794), .B1(r1[11]), .B2(n625), .C1(r1[10]), 
        .C2(n789), .ZN(n395) );
  AOI222_X1 U518 ( .A1(r1[8]), .A2(n788), .B1(r1[16]), .B2(n779), .C1(r1[15]), 
        .C2(n791), .ZN(n397) );
  NAND4_X1 U519 ( .A1(n327), .A2(n328), .A3(n329), .A4(n330), .ZN(N2069) );
  AOI222_X1 U520 ( .A1(n769), .A2(n730), .B1(n759), .B2(n723), .C1(n770), .C2(
        n715), .ZN(n330) );
  AOI21_X1 U521 ( .B1(r1[10]), .B2(n601), .A(n748), .ZN(n327) );
  AOI221_X1 U522 ( .B1(n755), .B2(n710), .C1(n767), .C2(n704), .A(n331), .ZN(
        n329) );
  AOI21_X1 U523 ( .B1(n440), .B2(n441), .A(n747), .ZN(n439) );
  AOI221_X1 U532 ( .B1(n755), .B2(r1[20]), .C1(n767), .C2(r1[19]), .A(n449), 
        .ZN(n440) );
  OAI222_X1 U541 ( .A1(n697), .A2(n319), .B1(n699), .B2(n366), .C1(n702), .C2(
        n332), .ZN(n449) );
  AOI22_X1 U542 ( .A1(n790), .A2(n683), .B1(n760), .B2(r1[19]), .ZN(n425) );
  AOI221_X1 U543 ( .B1(n755), .B2(n690), .C1(n767), .C2(r1[20]), .A(n428), 
        .ZN(n427) );
  AOI222_X1 U544 ( .A1(n770), .A2(n693), .B1(n214), .B2(n429), .C1(n759), .C2(
        n696), .ZN(n426) );
  INV_X1 U545 ( .A(r1[23]), .ZN(n697) );
  AOI222_X1 U546 ( .A1(n755), .A2(n715), .B1(n759), .B2(n729), .C1(n770), .C2(
        n725), .ZN(n315) );
  AOI211_X1 U547 ( .C1(r1[11]), .C2(n601), .A(n317), .B(n748), .ZN(n316) );
  AOI22_X1 U548 ( .A1(n767), .A2(n710), .B1(n320), .B2(n745), .ZN(n314) );
  BUF_X1 U549 ( .A(r1[17]), .Z(n680) );
  AOI22_X1 U550 ( .A1(n779), .A2(n736), .B1(n791), .B2(n728), .ZN(n179) );
  AOI22_X1 U551 ( .A1(n182), .A2(n118), .B1(n183), .B2(n157), .ZN(n180) );
  AOI221_X1 U552 ( .B1(n771), .B2(r1[27]), .C1(n762), .C2(n704), .A(n438), 
        .ZN(n437) );
  AOI21_X1 U553 ( .B1(r1[3]), .B2(n601), .A(n423), .ZN(n435) );
  BUF_X1 U554 ( .A(r1[17]), .Z(n681) );
  OAI21_X1 U555 ( .B1(n452), .B2(n453), .A(n766), .ZN(n450) );
  OAI221_X1 U556 ( .B1(n711), .B2(n386), .C1(n740), .C2(n455), .A(n456), .ZN(
        n453) );
  BUF_X1 U557 ( .A(r1[29]), .Z(n720) );
  BUF_X1 U558 ( .A(r1[29]), .Z(n721) );
  AOI22_X1 U559 ( .A1(n609), .A2(r1[20]), .B1(n624), .B2(n687), .ZN(n364) );
  AOI22_X1 U560 ( .A1(r1[15]), .A2(n781), .B1(r1[16]), .B2(n624), .ZN(n448) );
  AOI22_X1 U561 ( .A1(n677), .A2(n609), .B1(r1[15]), .B2(n624), .ZN(n467) );
  INV_X1 U562 ( .A(log), .ZN(n752) );
  NAND2_X1 U563 ( .A1(n499), .A2(n490), .ZN(n153) );
  OAI211_X1 U564 ( .C1(n101), .C2(n670), .A(n343), .B(n354), .ZN(N2067) );
  AOI22_X1 U565 ( .A1(n152), .A2(n642), .B1(n786), .B2(n728), .ZN(n151) );
  AOI222_X1 U566 ( .A1(n693), .A2(n574), .B1(n793), .B2(n698), .C1(n696), .C2(
        n786), .ZN(n241) );
  AOI222_X1 U567 ( .A1(r1[10]), .A2(n786), .B1(r1[11]), .B2(n793), .C1(r1[12]), 
        .C2(n787), .ZN(n431) );
  AOI222_X1 U568 ( .A1(n674), .A2(n786), .B1(n677), .B2(n793), .C1(r1[15]), 
        .C2(n787), .ZN(n379) );
  AOI222_X1 U569 ( .A1(r1[12]), .A2(n786), .B1(n674), .B2(n793), .C1(n678), 
        .C2(n787), .ZN(n396) );
  AOI22_X1 U570 ( .A1(n698), .A2(n786), .B1(n696), .B2(n574), .ZN(n235) );
  AOI22_X1 U571 ( .A1(n786), .A2(n700), .B1(n698), .B2(n574), .ZN(n220) );
  CLKBUF_X1 U572 ( .A(n197), .Z(n643) );
  NAND2_X1 U573 ( .A1(n478), .A2(n651), .ZN(n197) );
  OAI22_X1 U574 ( .A1(n195), .A2(n792), .B1(n196), .B2(n736), .ZN(n194) );
  OAI22_X1 U575 ( .A1(n726), .A2(n196), .B1(n792), .B2(n231), .ZN(n226) );
  AOI22_X1 U576 ( .A1(n733), .A2(n792), .B1(n196), .B2(n216), .ZN(n210) );
  OAI221_X1 U577 ( .B1(n654), .B2(n803), .C1(n695), .C2(n196), .A(n326), .ZN(
        n322) );
  OAI221_X1 U578 ( .B1(n682), .B2(n654), .C1(n711), .C2(n196), .A(n255), .ZN(
        n250) );
  OAI221_X1 U579 ( .B1(n654), .B2(n801), .C1(n702), .C2(n196), .A(n277), .ZN(
        n273) );
  OAI221_X1 U580 ( .B1(n654), .B2(n672), .C1(n802), .C2(n196), .A(n352), .ZN(
        n348) );
  AOI21_X1 U581 ( .B1(n196), .B2(n202), .A(n739), .ZN(n183) );
  OAI221_X1 U582 ( .B1(n654), .B2(n800), .C1(n709), .C2(n196), .A(n263), .ZN(
        n259) );
  OAI221_X1 U583 ( .B1(n654), .B2(n673), .C1(n691), .C2(n196), .A(n340), .ZN(
        n336) );
  OAI221_X1 U584 ( .B1(n654), .B2(n676), .C1(n697), .C2(n196), .A(n313), .ZN(
        n309) );
  OAI221_X1 U585 ( .B1(n573), .B2(n679), .C1(n699), .C2(n196), .A(n295), .ZN(
        n291) );
  AOI22_X1 U587 ( .A1(r1[1]), .A2(n600), .B1(r1[2]), .B2(n601), .ZN(n451) );
  OR3_X1 U588 ( .A1(n648), .A2(n600), .A3(n100), .ZN(n102) );
  AOI22_X1 U589 ( .A1(r1[0]), .A2(n600), .B1(r1[1]), .B2(n601), .ZN(n470) );
  AOI22_X1 U590 ( .A1(r1[26]), .A2(n600), .B1(r1[27]), .B2(n601), .ZN(n122) );
  AOI22_X1 U591 ( .A1(n246), .A2(n745), .B1(r1[15]), .B2(n600), .ZN(n245) );
  AOI22_X1 U592 ( .A1(n143), .A2(n746), .B1(n698), .B2(n600), .ZN(n142) );
  AOI22_X1 U593 ( .A1(n767), .A2(n727), .B1(n674), .B2(n600), .ZN(n265) );
  AOI22_X1 U594 ( .A1(n762), .A2(n727), .B1(r1[6]), .B2(n600), .ZN(n367) );
  AOI22_X1 U595 ( .A1(n134), .A2(n212), .B1(n684), .B2(n600), .ZN(n208) );
  AOI221_X1 U596 ( .B1(r1[20]), .B2(n600), .C1(n689), .C2(n601), .A(n116), 
        .ZN(n181) );
  AOI221_X1 U597 ( .B1(r1[2]), .B2(n600), .C1(n772), .C2(n776), .A(n439), .ZN(
        n436) );
  AOI222_X1 U598 ( .A1(n677), .A2(n600), .B1(n745), .B2(n257), .C1(n767), .C2(
        n736), .ZN(n256) );
  AOI222_X1 U599 ( .A1(r1[16]), .A2(n600), .B1(n229), .B2(n238), .C1(n790), 
        .C2(n776), .ZN(n237) );
  AOI221_X1 U600 ( .B1(n688), .B2(n600), .C1(n694), .C2(n601), .A(n116), .ZN(
        n170) );
  AOI221_X1 U601 ( .B1(n710), .B2(n600), .C1(r1[28]), .C2(n601), .A(n116), 
        .ZN(n115) );
  AOI221_X1 U602 ( .B1(n696), .B2(n600), .C1(n793), .C2(n776), .A(n149), .ZN(
        n148) );
  AOI222_X1 U603 ( .A1(n704), .A2(n601), .B1(n134), .B2(n579), .C1(r1[25]), 
        .C2(n600), .ZN(n133) );
  NOR4_X1 U604 ( .A1(n297), .A2(n648), .A3(n601), .A4(n600), .ZN(n128) );
  BUF_X1 U605 ( .A(n99), .Z(n647) );
  AOI22_X1 U606 ( .A1(n111), .A2(n107), .B1(n112), .B2(n784), .ZN(n109) );
  AND4_X1 U607 ( .A1(n105), .A2(n761), .A3(n106), .A4(n107), .ZN(n104) );
  AOI22_X1 U608 ( .A1(n693), .A2(n107), .B1(n696), .B2(n788), .ZN(n188) );
  AOI22_X1 U609 ( .A1(r1[26]), .A2(n107), .B1(n786), .B2(n736), .ZN(n146) );
  AOI221_X1 U610 ( .B1(n696), .B2(n107), .C1(n698), .C2(n788), .A(n175), .ZN(
        n173) );
  INV_X1 U611 ( .A(n107), .ZN(n784) );
  AOI22_X1 U612 ( .A1(n689), .A2(n107), .B1(n786), .B2(n704), .ZN(n203) );
  CLKBUF_X1 U613 ( .A(n168), .Z(n645) );
  NAND2_X1 U614 ( .A1(n478), .A2(n653), .ZN(n168) );
  NAND2_X1 U615 ( .A1(n478), .A2(n481), .ZN(n408) );
  NAND2_X1 U616 ( .A1(n481), .A2(n491), .ZN(n287) );
  NAND2_X1 U617 ( .A1(n481), .A2(n499), .ZN(n332) );
  NAND2_X1 U618 ( .A1(n481), .A2(n497), .ZN(n319) );
  NAND2_X1 U619 ( .A1(n482), .A2(n481), .ZN(n476) );
  OAI22_X1 U620 ( .A1(n733), .A2(n607), .B1(n722), .B2(n640), .ZN(n175) );
  OAI222_X1 U621 ( .A1(n607), .A2(n799), .B1(n640), .B2(n685), .C1(n642), .C2(
        n682), .ZN(n324) );
  OAI222_X1 U622 ( .A1(n699), .A2(n607), .B1(n640), .B2(n697), .C1(n642), .C2(
        n695), .ZN(n252) );
  OAI222_X1 U623 ( .A1(n607), .A2(n695), .B1(n640), .B2(n691), .C1(n642), .C2(
        n802), .ZN(n275) );
  OAI222_X1 U624 ( .A1(n607), .A2(n682), .B1(n640), .B2(n800), .C1(n642), .C2(
        n801), .ZN(n350) );
  OAI222_X1 U625 ( .A1(n697), .A2(n607), .B1(n640), .B2(n695), .C1(n642), .C2(
        n691), .ZN(n261) );
  OAI222_X1 U626 ( .A1(n607), .A2(n685), .B1(n640), .B2(n682), .C1(n642), .C2(
        n800), .ZN(n338) );
  OAI222_X1 U627 ( .A1(n607), .A2(n672), .B1(n640), .B2(n671), .C1(n642), .C2(
        n670), .ZN(n465) );
  OAI221_X1 U628 ( .B1(n702), .B2(n640), .C1(n709), .C2(n607), .A(n235), .ZN(
        n234) );
  OAI222_X1 U629 ( .A1(n607), .A2(n671), .B1(n640), .B2(n670), .C1(n642), .C2(
        n669), .ZN(n494) );
  OAI222_X1 U630 ( .A1(n607), .A2(n676), .B1(n640), .B2(n803), .C1(n642), .C2(
        n673), .ZN(n415) );
  OAI221_X1 U631 ( .B1(n705), .B2(n640), .C1(n714), .C2(n607), .A(n220), .ZN(
        n219) );
  OAI222_X1 U632 ( .A1(n607), .A2(n673), .B1(n640), .B2(n672), .C1(n642), .C2(
        n671), .ZN(n446) );
  OAI222_X1 U633 ( .A1(n607), .A2(n802), .B1(n640), .B2(n799), .C1(n642), .C2(
        n685), .ZN(n311) );
  OAI222_X1 U634 ( .A1(n607), .A2(n800), .B1(n640), .B2(n801), .C1(n642), .C2(
        n679), .ZN(n362) );
  OAI222_X1 U635 ( .A1(n607), .A2(n691), .B1(n640), .B2(n802), .C1(n642), .C2(
        n799), .ZN(n293) );
  INV_X1 U636 ( .A(n177), .ZN(n793) );
  NAND2_X1 U637 ( .A1(n176), .A2(n177), .ZN(n150) );
  NAND4_X1 U638 ( .A1(n504), .A2(n501), .A3(n503), .A4(n502), .ZN(n99) );
  AND4_X2 U639 ( .A1(n136), .A2(n108), .A3(n137), .A4(n138), .ZN(n107) );
  INV_X1 U640 ( .A(n626), .ZN(n785) );
  NAND2_X1 U641 ( .A1(n489), .A2(n606), .ZN(n108) );
  NAND2_X1 U642 ( .A1(n497), .A2(n651), .ZN(n137) );
  NAND2_X1 U643 ( .A1(n497), .A2(n652), .ZN(n138) );
  AOI22_X1 U644 ( .A1(n574), .A2(n776), .B1(n112), .B2(n785), .ZN(n132) );
  NAND2_X1 U645 ( .A1(n737), .A2(n785), .ZN(n129) );
  NOR3_X1 U646 ( .A1(n119), .A2(n789), .A3(n785), .ZN(n113) );
  AOI221_X1 U647 ( .B1(r1[8]), .B2(n778), .C1(n683), .C2(n792), .A(n382), .ZN(
        n381) );
  INV_X1 U648 ( .A(n573), .ZN(n778) );
  NOR3_X1 U649 ( .A1(n786), .A2(n625), .A3(n150), .ZN(n136) );
  AOI211_X1 U650 ( .C1(n128), .C2(n279), .A(n162), .B(n280), .ZN(n278) );
  INV_X1 U651 ( .A(r2[0]), .ZN(n798) );
  OAI21_X1 U652 ( .B1(n389), .B2(n390), .A(n391), .ZN(n388) );
  INV_X1 U653 ( .A(r1[2]), .ZN(n664) );
  INV_X1 U654 ( .A(r1[3]), .ZN(n665) );
  INV_X1 U655 ( .A(r1[4]), .ZN(n666) );
  INV_X1 U656 ( .A(r1[5]), .ZN(n667) );
  INV_X1 U657 ( .A(r1[6]), .ZN(n668) );
  INV_X1 U658 ( .A(r1[7]), .ZN(n669) );
  INV_X1 U659 ( .A(r1[8]), .ZN(n670) );
  INV_X1 U660 ( .A(r1[9]), .ZN(n671) );
  INV_X1 U661 ( .A(r1[10]), .ZN(n672) );
  INV_X1 U662 ( .A(r1[11]), .ZN(n673) );
  CLKBUF_X1 U663 ( .A(r1[21]), .Z(n686) );
  CLKBUF_X1 U664 ( .A(r1[21]), .Z(n687) );
  CLKBUF_X1 U665 ( .A(r1[21]), .Z(n688) );
  CLKBUF_X1 U666 ( .A(r1[21]), .Z(n689) );
  CLKBUF_X1 U667 ( .A(r1[21]), .Z(n690) );
  INV_X1 U668 ( .A(n697), .ZN(n696) );
  INV_X1 U669 ( .A(n699), .ZN(n698) );
  INV_X1 U670 ( .A(r1[25]), .ZN(n701) );
  INV_X1 U671 ( .A(r1[25]), .ZN(n702) );
  INV_X1 U672 ( .A(r1[25]), .ZN(n703) );
  INV_X1 U673 ( .A(r1[26]), .ZN(n705) );
  INV_X1 U674 ( .A(r1[26]), .ZN(n706) );
  INV_X1 U675 ( .A(r1[26]), .ZN(n707) );
  INV_X1 U676 ( .A(r1[26]), .ZN(n708) );
  INV_X1 U677 ( .A(r1[26]), .ZN(n709) );
  INV_X1 U678 ( .A(r1[27]), .ZN(n711) );
  INV_X1 U679 ( .A(r1[27]), .ZN(n712) );
  INV_X1 U680 ( .A(r1[27]), .ZN(n713) );
  INV_X1 U681 ( .A(r1[27]), .ZN(n714) );
  INV_X1 U682 ( .A(r1[28]), .ZN(n716) );
  INV_X1 U683 ( .A(r1[28]), .ZN(n717) );
  INV_X1 U684 ( .A(r1[28]), .ZN(n718) );
  INV_X1 U685 ( .A(r1[28]), .ZN(n719) );
  CLKBUF_X1 U686 ( .A(r1[31]), .Z(n734) );
  CLKBUF_X1 U687 ( .A(r1[31]), .Z(n735) );
  INV_X1 U688 ( .A(n741), .ZN(n737) );
  INV_X1 U689 ( .A(n734), .ZN(n738) );
  INV_X1 U690 ( .A(n735), .ZN(n739) );
  INV_X1 U691 ( .A(n735), .ZN(n740) );
  INV_X1 U692 ( .A(r1[31]), .ZN(n741) );
  INV_X2 U693 ( .A(n270), .ZN(n755) );
  INV_X2 U694 ( .A(n287), .ZN(n767) );
  INV_X2 U695 ( .A(n153), .ZN(n786) );
endmodule


module comparator_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n202, n292, n65, n66, n69, n71, n72, n74, n75, n77, n80, n81, n83,
         n84, n86, n87, n89, n92, n93, n95, n96, n98, n99, n101, n104, n105,
         n108, n110, n111, n113, n116, n117, n120, n122, n123, n125, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, net52631, net52642,
         net52646, net52650, net52651, net52652, net54692, n203, n204, n205,
         n206, n207, n208, n209, n210, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291;

  XOR2_X1 U101 ( .A(A[30]), .B(net52651), .Z(n69) );
  NAND3_X1 U170 ( .A1(n196), .A2(n149), .A3(n146), .ZN(n195) );
  NAND3_X1 U174 ( .A1(n199), .A2(n198), .A3(n283), .ZN(n196) );
  AND2_X1 U1 ( .A1(n89), .A2(n92), .ZN(n226) );
  NAND2_X1 U2 ( .A1(n86), .A2(n207), .ZN(n228) );
  NOR2_X1 U3 ( .A1(n84), .A2(n81), .ZN(n244) );
  NAND2_X1 U4 ( .A1(n83), .A2(n243), .ZN(n242) );
  INV_X1 U5 ( .A(n87), .ZN(n243) );
  NAND2_X1 U6 ( .A1(n125), .A2(n128), .ZN(n216) );
  OAI21_X1 U7 ( .B1(n215), .B2(n234), .A(n235), .ZN(n219) );
  NOR2_X1 U8 ( .A1(n123), .A2(n208), .ZN(n235) );
  NAND2_X1 U9 ( .A1(n122), .A2(n203), .ZN(n234) );
  NOR2_X1 U10 ( .A1(n210), .A2(n216), .ZN(n215) );
  NOR2_X1 U11 ( .A1(n120), .A2(n117), .ZN(n218) );
  NAND2_X1 U12 ( .A1(n113), .A2(n116), .ZN(n220) );
  OAI21_X1 U13 ( .B1(n217), .B2(n236), .A(n237), .ZN(n248) );
  NOR2_X1 U14 ( .A1(n111), .A2(n209), .ZN(n237) );
  NAND2_X1 U15 ( .A1(n110), .A2(n205), .ZN(n236) );
  AOI21_X1 U16 ( .B1(n218), .B2(n219), .A(n220), .ZN(n217) );
  NOR2_X1 U17 ( .A1(n108), .A2(n105), .ZN(n238) );
  AOI21_X1 U18 ( .B1(n222), .B2(n223), .A(n224), .ZN(n221) );
  AND2_X1 U19 ( .A1(n101), .A2(n104), .ZN(n222) );
  NAND2_X1 U20 ( .A1(n98), .A2(n206), .ZN(n224) );
  NAND2_X1 U21 ( .A1(n238), .A2(n248), .ZN(n223) );
  NOR2_X1 U22 ( .A1(n96), .A2(n93), .ZN(n241) );
  NAND2_X1 U23 ( .A1(n95), .A2(n240), .ZN(n239) );
  INV_X1 U24 ( .A(n99), .ZN(n240) );
  AND2_X1 U25 ( .A1(n77), .A2(n80), .ZN(n230) );
  NAND2_X1 U26 ( .A1(n74), .A2(n204), .ZN(n232) );
  NOR2_X1 U27 ( .A1(n72), .A2(n233), .ZN(n247) );
  INV_X1 U28 ( .A(n69), .ZN(n233) );
  NAND2_X1 U29 ( .A1(n71), .A2(n246), .ZN(n245) );
  INV_X1 U30 ( .A(n75), .ZN(n246) );
  OR2_X1 U31 ( .A1(n262), .A2(B[11]), .ZN(n203) );
  OR2_X1 U32 ( .A1(n273), .A2(B[27]), .ZN(n204) );
  OR2_X1 U33 ( .A1(n289), .A2(B[15]), .ZN(n205) );
  OR2_X1 U34 ( .A1(n287), .A2(B[19]), .ZN(n206) );
  OR2_X1 U35 ( .A1(n269), .A2(B[23]), .ZN(n207) );
  AND2_X1 U36 ( .A1(B[13]), .A2(n263), .ZN(n208) );
  AND2_X1 U37 ( .A1(B[17]), .A2(n265), .ZN(n209) );
  AND2_X1 U38 ( .A1(n127), .A2(net52631), .ZN(n210) );
  CLKBUF_X1 U39 ( .A(n276), .Z(LE) );
  AOI21_X1 U40 ( .B1(n230), .B2(n231), .A(n232), .ZN(n229) );
  OAI21_X1 U41 ( .B1(n225), .B2(n242), .A(n244), .ZN(n231) );
  NAND2_X1 U42 ( .A1(n213), .A2(n214), .ZN(net52652) );
  AOI21_X1 U43 ( .B1(n226), .B2(n227), .A(n228), .ZN(n225) );
  NOR2_X1 U44 ( .A1(n252), .A2(B[0]), .ZN(n212) );
  OAI21_X1 U45 ( .B1(n229), .B2(n245), .A(n247), .ZN(n214) );
  OAI21_X1 U46 ( .B1(n221), .B2(n239), .A(n241), .ZN(n227) );
  NAND2_X1 U47 ( .A1(B[30]), .A2(net54692), .ZN(n213) );
  OR2_X1 U48 ( .A1(B[2]), .A2(n253), .ZN(n198) );
  AOI21_X1 U49 ( .B1(net52652), .B2(n65), .A(n66), .ZN(GE) );
  NAND2_X1 U50 ( .A1(B[0]), .A2(n250), .ZN(n154) );
  AND2_X1 U51 ( .A1(n252), .A2(n251), .ZN(n250) );
  INV_X1 U52 ( .A(A[1]), .ZN(n251) );
  NOR2_X1 U53 ( .A1(n192), .A2(n135), .ZN(n134) );
  NOR2_X1 U54 ( .A1(n192), .A2(n132), .ZN(n188) );
  INV_X1 U55 ( .A(n95), .ZN(net52642) );
  INV_X1 U56 ( .A(n131), .ZN(n278) );
  INV_X1 U57 ( .A(n141), .ZN(n281) );
  INV_X1 U58 ( .A(n129), .ZN(net52631) );
  OAI211_X1 U59 ( .C1(n166), .C2(n167), .A(n89), .B(n86), .ZN(n165) );
  NAND2_X1 U60 ( .A1(n207), .A2(n169), .ZN(n167) );
  AOI211_X1 U61 ( .C1(n171), .C2(n170), .A(n93), .B(net52642), .ZN(n166) );
  OAI211_X1 U62 ( .C1(n160), .C2(n161), .A(n77), .B(n74), .ZN(n159) );
  NAND2_X1 U63 ( .A1(n204), .A2(n163), .ZN(n161) );
  AOI211_X1 U64 ( .C1(n165), .C2(n164), .A(n81), .B(net52646), .ZN(n160) );
  OAI211_X1 U65 ( .C1(n178), .C2(n179), .A(n113), .B(n110), .ZN(n177) );
  NAND2_X1 U66 ( .A1(n205), .A2(n181), .ZN(n179) );
  AOI211_X1 U67 ( .C1(n183), .C2(n182), .A(n117), .B(n208), .ZN(n178) );
  OAI211_X1 U68 ( .C1(n184), .C2(n185), .A(n125), .B(n122), .ZN(n183) );
  NAND2_X1 U69 ( .A1(n203), .A2(n187), .ZN(n185) );
  AOI211_X1 U70 ( .C1(n189), .C2(n188), .A(n129), .B(n278), .ZN(n184) );
  NOR2_X1 U71 ( .A1(n260), .A2(B[9]), .ZN(n132) );
  OAI211_X1 U72 ( .C1(n172), .C2(n173), .A(n101), .B(n98), .ZN(n171) );
  NAND2_X1 U73 ( .A1(n206), .A2(n175), .ZN(n173) );
  AOI211_X1 U74 ( .C1(n177), .C2(n176), .A(n105), .B(n209), .ZN(n172) );
  NOR2_X1 U75 ( .A1(n162), .A2(n75), .ZN(n74) );
  NOR2_X1 U76 ( .A1(n186), .A2(n123), .ZN(n122) );
  NOR2_X1 U77 ( .A1(n180), .A2(n111), .ZN(n110) );
  NOR2_X1 U78 ( .A1(n174), .A2(n99), .ZN(n98) );
  NOR2_X1 U79 ( .A1(n168), .A2(n87), .ZN(n86) );
  NAND2_X1 U80 ( .A1(B[9]), .A2(n260), .ZN(n131) );
  NOR2_X1 U81 ( .A1(n197), .A2(n147), .ZN(n146) );
  NOR2_X1 U82 ( .A1(n162), .A2(n72), .ZN(n158) );
  NOR2_X1 U83 ( .A1(n197), .A2(n144), .ZN(n194) );
  NOR2_X1 U84 ( .A1(n186), .A2(n120), .ZN(n182) );
  NOR2_X1 U85 ( .A1(n180), .A2(n108), .ZN(n176) );
  NOR2_X1 U86 ( .A1(n174), .A2(n96), .ZN(n170) );
  NOR2_X1 U87 ( .A1(n168), .A2(n84), .ZN(n164) );
  NAND2_X1 U88 ( .A1(n169), .A2(n92), .ZN(n93) );
  NAND2_X1 U89 ( .A1(n163), .A2(n80), .ZN(n81) );
  NAND2_X1 U90 ( .A1(n193), .A2(n140), .ZN(n141) );
  NAND2_X1 U91 ( .A1(n187), .A2(n128), .ZN(n129) );
  NAND2_X1 U92 ( .A1(n175), .A2(n104), .ZN(n105) );
  NAND2_X1 U93 ( .A1(n181), .A2(n116), .ZN(n117) );
  AND2_X1 U94 ( .A1(n198), .A2(n153), .ZN(n152) );
  INV_X1 U95 ( .A(n143), .ZN(n282) );
  INV_X1 U96 ( .A(n83), .ZN(net52646) );
  INV_X1 U97 ( .A(n140), .ZN(n280) );
  INV_X1 U98 ( .A(n153), .ZN(n284) );
  NOR2_X1 U99 ( .A1(n255), .A2(B[4]), .ZN(n197) );
  NOR2_X1 U100 ( .A1(n288), .A2(B[16]), .ZN(n180) );
  NOR2_X1 U102 ( .A1(n270), .A2(B[24]), .ZN(n168) );
  NOR2_X1 U103 ( .A1(n291), .A2(B[12]), .ZN(n186) );
  NOR2_X1 U104 ( .A1(n290), .A2(B[20]), .ZN(n174) );
  NOR2_X1 U105 ( .A1(n275), .A2(B[29]), .ZN(n72) );
  NOR2_X1 U106 ( .A1(n254), .A2(B[3]), .ZN(n150) );
  OAI211_X1 U107 ( .C1(n190), .C2(n191), .A(n137), .B(n134), .ZN(n189) );
  NAND2_X1 U108 ( .A1(n279), .A2(n193), .ZN(n191) );
  AOI211_X1 U109 ( .C1(n194), .C2(n195), .A(n141), .B(n282), .ZN(n190) );
  INV_X1 U110 ( .A(n138), .ZN(n279) );
  NOR2_X1 U111 ( .A1(n256), .A2(B[5]), .ZN(n144) );
  NAND2_X1 U112 ( .A1(B[3]), .A2(n254), .ZN(n149) );
  NOR2_X1 U113 ( .A1(n258), .A2(B[7]), .ZN(n138) );
  NOR2_X1 U114 ( .A1(n265), .A2(B[17]), .ZN(n108) );
  NOR2_X1 U115 ( .A1(n271), .A2(B[25]), .ZN(n84) );
  NAND2_X1 U116 ( .A1(B[6]), .A2(n257), .ZN(n140) );
  NAND2_X1 U117 ( .A1(B[26]), .A2(n272), .ZN(n80) );
  NAND2_X1 U118 ( .A1(B[19]), .A2(n287), .ZN(n101) );
  NAND2_X1 U119 ( .A1(B[29]), .A2(n275), .ZN(n71) );
  OAI21_X1 U120 ( .B1(n156), .B2(n66), .A(n65), .ZN(n202) );
  AOI22_X1 U121 ( .A1(A[30]), .A2(net52651), .B1(n157), .B2(n69), .ZN(n156) );
  AOI21_X1 U122 ( .B1(n159), .B2(n158), .A(net52650), .ZN(n157) );
  INV_X1 U123 ( .A(n71), .ZN(net52650) );
  NAND2_X1 U124 ( .A1(B[11]), .A2(n262), .ZN(n125) );
  NAND2_X1 U125 ( .A1(B[10]), .A2(n261), .ZN(n128) );
  NAND2_X1 U126 ( .A1(B[18]), .A2(n266), .ZN(n104) );
  NAND2_X1 U127 ( .A1(B[14]), .A2(n264), .ZN(n116) );
  NAND2_X1 U128 ( .A1(B[5]), .A2(n256), .ZN(n143) );
  NAND2_X1 U129 ( .A1(B[7]), .A2(n258), .ZN(n137) );
  NAND2_X1 U130 ( .A1(B[27]), .A2(n273), .ZN(n77) );
  NAND2_X1 U131 ( .A1(B[23]), .A2(n269), .ZN(n89) );
  NAND2_X1 U132 ( .A1(B[25]), .A2(n271), .ZN(n83) );
  NAND2_X1 U133 ( .A1(B[15]), .A2(n289), .ZN(n113) );
  OR2_X1 U134 ( .A1(n272), .A2(B[26]), .ZN(n163) );
  OR2_X1 U135 ( .A1(n257), .A2(B[6]), .ZN(n193) );
  NAND2_X1 U136 ( .A1(B[2]), .A2(n253), .ZN(n153) );
  INV_X1 U137 ( .A(B[31]), .ZN(n277) );
  AND2_X1 U138 ( .A1(B[4]), .A2(n255), .ZN(n147) );
  OR2_X1 U139 ( .A1(n261), .A2(B[10]), .ZN(n187) );
  OR2_X1 U140 ( .A1(n266), .A2(B[18]), .ZN(n175) );
  OR2_X1 U141 ( .A1(n264), .A2(B[14]), .ZN(n181) );
  AND2_X1 U142 ( .A1(B[12]), .A2(n291), .ZN(n123) );
  AND2_X1 U143 ( .A1(B[16]), .A2(n288), .ZN(n111) );
  INV_X1 U144 ( .A(B[30]), .ZN(net52651) );
  AND2_X1 U145 ( .A1(B[20]), .A2(n290), .ZN(n99) );
  AND2_X1 U146 ( .A1(B[24]), .A2(n270), .ZN(n87) );
  INV_X1 U147 ( .A(B[1]), .ZN(n286) );
  INV_X1 U148 ( .A(n202), .ZN(n276) );
  INV_X1 U149 ( .A(A[19]), .ZN(n287) );
  NOR2_X1 U150 ( .A1(n277), .A2(A[31]), .ZN(n66) );
  INV_X1 U151 ( .A(A[16]), .ZN(n288) );
  INV_X1 U152 ( .A(A[15]), .ZN(n289) );
  INV_X1 U153 ( .A(A[12]), .ZN(n291) );
  INV_X1 U154 ( .A(A[20]), .ZN(n290) );
  NAND2_X1 U155 ( .A1(A[31]), .A2(n277), .ZN(n65) );
  INV_X1 U156 ( .A(n150), .ZN(n283) );
  OAI211_X1 U157 ( .C1(A[1]), .C2(n212), .A(n285), .B(n152), .ZN(n199) );
  INV_X1 U158 ( .A(n201), .ZN(n285) );
  AOI21_X1 U159 ( .B1(n200), .B2(A[1]), .A(n286), .ZN(n201) );
  AOI21_X1 U160 ( .B1(net52652), .B2(n65), .A(n66), .ZN(n292) );
  NOR2_X1 U161 ( .A1(n263), .A2(B[13]), .ZN(n120) );
  AOI21_X1 U162 ( .B1(n152), .B2(n151), .A(n284), .ZN(n148) );
  AOI22_X1 U163 ( .A1(n286), .A2(n154), .B1(n155), .B2(A[1]), .ZN(n151) );
  AOI21_X1 U164 ( .B1(n130), .B2(n131), .A(n132), .ZN(n127) );
  AOI21_X1 U165 ( .B1(n133), .B2(n134), .A(n135), .ZN(n130) );
  AOI21_X1 U166 ( .B1(n136), .B2(n137), .A(n138), .ZN(n133) );
  OR2_X1 U167 ( .A1(n268), .A2(B[22]), .ZN(n169) );
  NAND2_X1 U168 ( .A1(B[22]), .A2(n268), .ZN(n92) );
  NOR2_X1 U169 ( .A1(n274), .A2(B[28]), .ZN(n162) );
  AND2_X1 U171 ( .A1(B[28]), .A2(n274), .ZN(n75) );
  AOI21_X1 U172 ( .B1(n142), .B2(n143), .A(n144), .ZN(n139) );
  AOI21_X1 U173 ( .B1(n148), .B2(n149), .A(n150), .ZN(n145) );
  NAND2_X1 U175 ( .A1(B[21]), .A2(n267), .ZN(n95) );
  NOR2_X1 U176 ( .A1(n267), .A2(B[21]), .ZN(n96) );
  AND2_X1 U177 ( .A1(n292), .A2(n276), .ZN(EQ) );
  AOI21_X1 U178 ( .B1(n139), .B2(n281), .A(n280), .ZN(n136) );
  NOR2_X1 U179 ( .A1(n252), .A2(B[0]), .ZN(n200) );
  AOI21_X1 U180 ( .B1(n145), .B2(n146), .A(n147), .ZN(n142) );
  NAND2_X1 U181 ( .A1(B[0]), .A2(n252), .ZN(n155) );
  NOR2_X1 U182 ( .A1(n259), .A2(B[8]), .ZN(n192) );
  AND2_X1 U183 ( .A1(B[8]), .A2(n259), .ZN(n135) );
  INV_X1 U184 ( .A(A[0]), .ZN(n252) );
  INV_X1 U185 ( .A(A[2]), .ZN(n253) );
  INV_X1 U186 ( .A(A[3]), .ZN(n254) );
  INV_X1 U187 ( .A(A[4]), .ZN(n255) );
  INV_X1 U188 ( .A(A[5]), .ZN(n256) );
  INV_X1 U189 ( .A(A[6]), .ZN(n257) );
  INV_X1 U190 ( .A(A[7]), .ZN(n258) );
  INV_X1 U191 ( .A(A[8]), .ZN(n259) );
  INV_X1 U192 ( .A(A[9]), .ZN(n260) );
  INV_X1 U193 ( .A(A[10]), .ZN(n261) );
  INV_X1 U194 ( .A(A[11]), .ZN(n262) );
  INV_X1 U195 ( .A(A[13]), .ZN(n263) );
  INV_X1 U196 ( .A(A[14]), .ZN(n264) );
  INV_X1 U197 ( .A(A[17]), .ZN(n265) );
  INV_X1 U198 ( .A(A[18]), .ZN(n266) );
  INV_X1 U199 ( .A(A[21]), .ZN(n267) );
  INV_X1 U200 ( .A(A[22]), .ZN(n268) );
  INV_X1 U201 ( .A(A[23]), .ZN(n269) );
  INV_X1 U202 ( .A(A[24]), .ZN(n270) );
  INV_X1 U203 ( .A(A[25]), .ZN(n271) );
  INV_X1 U204 ( .A(A[26]), .ZN(n272) );
  INV_X1 U205 ( .A(A[27]), .ZN(n273) );
  INV_X1 U206 ( .A(A[28]), .ZN(n274) );
  INV_X1 U207 ( .A(A[29]), .ZN(n275) );
  INV_X1 U208 ( .A(A[30]), .ZN(net54692) );
endmodule


module comparator ( r1, r2, sel, data_out );
  input [31:0] r1;
  input [31:0] r2;
  input [2:0] sel;
  output [31:0] data_out;
  wire   N26, N27, N28, n5, n6, n8, net52585, n7, n9, n10, n11, n12, n13;
  assign data_out[31] = 1'b0;
  assign data_out[30] = 1'b0;
  assign data_out[29] = 1'b0;
  assign data_out[28] = 1'b0;
  assign data_out[27] = 1'b0;
  assign data_out[26] = 1'b0;
  assign data_out[25] = 1'b0;
  assign data_out[24] = 1'b0;
  assign data_out[23] = 1'b0;
  assign data_out[22] = 1'b0;
  assign data_out[21] = 1'b0;
  assign data_out[20] = 1'b0;
  assign data_out[19] = 1'b0;
  assign data_out[18] = 1'b0;
  assign data_out[17] = 1'b0;
  assign data_out[16] = 1'b0;
  assign data_out[15] = 1'b0;
  assign data_out[14] = 1'b0;
  assign data_out[13] = 1'b0;
  assign data_out[12] = 1'b0;
  assign data_out[11] = 1'b0;
  assign data_out[10] = 1'b0;
  assign data_out[9] = 1'b0;
  assign data_out[8] = 1'b0;
  assign data_out[7] = 1'b0;
  assign data_out[6] = 1'b0;
  assign data_out[5] = 1'b0;
  assign data_out[4] = 1'b0;
  assign data_out[3] = 1'b0;
  assign data_out[2] = 1'b0;
  assign data_out[1] = 1'b0;

  comparator_DW01_cmp6_0 r69 ( .A(r1), .B(r2), .TC(1'b0), .EQ(N26), .LE(N27), 
        .GE(N28) );
  NAND2_X1 U2 ( .A1(N26), .A2(n7), .ZN(n9) );
  NAND2_X1 U4 ( .A1(N27), .A2(sel[0]), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(net52585) );
  INV_X1 U6 ( .A(sel[0]), .ZN(n7) );
  OR2_X1 U7 ( .A1(n12), .A2(n11), .ZN(n6) );
  NAND2_X1 U8 ( .A1(sel[2]), .A2(n13), .ZN(n11) );
  XNOR2_X1 U9 ( .A(N28), .B(n7), .ZN(n8) );
  MUX2_X1 U10 ( .A(N27), .B(N26), .S(n7), .Z(n12) );
  AOI22_X1 U11 ( .A1(sel[1]), .A2(n8), .B1(net52585), .B2(n13), .ZN(n5) );
  INV_X1 U12 ( .A(sel[1]), .ZN(n13) );
  OAI21_X1 U13 ( .B1(n5), .B2(sel[2]), .A(n6), .ZN(data_out[0]) );
endmodule


module mux11to1_nbit32 ( A, B, C, D, E, F, H, sel, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [31:0] H;
  input [3:0] sel;
  output [31:0] Y;
  wire   n4, n5, n6, n7, n8, n9, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n107, n108, net52587, net56040, net56038, net56036, net56046,
         net56044, net56042, net56052, net56050, net56048, net56058, net56056,
         net56054, net56064, net56062, net56060, net56070, net56068, net56066,
         net56076, net56074, net56072, n11, n105, n10, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153;

  NAND3_X1 U110 ( .A1(n4), .A2(n5), .A3(n6), .ZN(Y[9]) );
  NAND3_X1 U111 ( .A1(n14), .A2(n15), .A3(n16), .ZN(Y[8]) );
  NAND3_X1 U113 ( .A1(n20), .A2(n21), .A3(n22), .ZN(Y[6]) );
  NAND3_X1 U115 ( .A1(n26), .A2(n27), .A3(n28), .ZN(Y[4]) );
  NAND3_X1 U116 ( .A1(n29), .A2(n30), .A3(n31), .ZN(Y[3]) );
  NAND3_X1 U118 ( .A1(n35), .A2(n36), .A3(n37), .ZN(Y[30]) );
  NAND3_X1 U119 ( .A1(n40), .A2(n39), .A3(n38), .ZN(Y[2]) );
  NAND3_X1 U120 ( .A1(n41), .A2(n42), .A3(n43), .ZN(Y[29]) );
  NAND3_X1 U121 ( .A1(n44), .A2(n45), .A3(n46), .ZN(Y[28]) );
  NAND3_X1 U122 ( .A1(n47), .A2(n48), .A3(n49), .ZN(Y[27]) );
  NAND3_X1 U123 ( .A1(n50), .A2(n51), .A3(n52), .ZN(Y[26]) );
  NAND3_X1 U124 ( .A1(n53), .A2(n54), .A3(n55), .ZN(Y[25]) );
  NAND3_X1 U125 ( .A1(n56), .A2(n57), .A3(n58), .ZN(Y[24]) );
  NAND3_X1 U126 ( .A1(n59), .A2(n60), .A3(n61), .ZN(Y[23]) );
  NAND3_X1 U127 ( .A1(n62), .A2(n63), .A3(n64), .ZN(Y[22]) );
  NAND3_X1 U128 ( .A1(n65), .A2(n66), .A3(n67), .ZN(Y[21]) );
  NAND3_X1 U129 ( .A1(n68), .A2(n69), .A3(n70), .ZN(Y[20]) );
  NAND3_X1 U130 ( .A1(n71), .A2(n72), .A3(n73), .ZN(Y[1]) );
  NAND3_X1 U131 ( .A1(n74), .A2(n75), .A3(n76), .ZN(Y[19]) );
  NAND3_X1 U132 ( .A1(n77), .A2(n78), .A3(n79), .ZN(Y[18]) );
  NAND3_X1 U133 ( .A1(n82), .A2(n81), .A3(n80), .ZN(Y[17]) );
  NAND3_X1 U134 ( .A1(n83), .A2(n84), .A3(n85), .ZN(Y[16]) );
  NAND3_X1 U135 ( .A1(n86), .A2(n87), .A3(n88), .ZN(Y[15]) );
  NAND3_X1 U136 ( .A1(n89), .A2(n90), .A3(n91), .ZN(Y[14]) );
  NAND3_X1 U137 ( .A1(n92), .A2(n93), .A3(n94), .ZN(Y[13]) );
  NAND3_X1 U140 ( .A1(n101), .A2(n102), .A3(n103), .ZN(Y[10]) );
  BUF_X1 U2 ( .A(n9), .Z(net56048) );
  BUF_X1 U3 ( .A(n9), .Z(net56050) );
  AND2_X1 U4 ( .A1(n131), .A2(n132), .ZN(n126) );
  AND2_X1 U5 ( .A1(n34), .A2(n33), .ZN(n109) );
  AND2_X1 U6 ( .A1(n95), .A2(n96), .ZN(n110) );
  AND2_X1 U7 ( .A1(n98), .A2(n99), .ZN(n111) );
  AND2_X1 U8 ( .A1(n17), .A2(n18), .ZN(n112) );
  INV_X1 U9 ( .A(n104), .ZN(n115) );
  AND2_X1 U10 ( .A1(n23), .A2(n24), .ZN(n113) );
  NOR2_X1 U11 ( .A1(n116), .A2(n115), .ZN(n114) );
  NAND3_X1 U12 ( .A1(n140), .A2(n141), .A3(n142), .ZN(n116) );
  AOI22_X1 U13 ( .A1(E[4]), .A2(net56070), .B1(C[4]), .B2(net56076), .ZN(n26)
         );
  NAND2_X1 U14 ( .A1(A[18]), .A2(net56036), .ZN(n117) );
  NAND2_X1 U15 ( .A1(B[18]), .A2(net56042), .ZN(n118) );
  NAND2_X1 U16 ( .A1(F[18]), .A2(net56048), .ZN(n119) );
  AND3_X1 U17 ( .A1(n117), .A2(n118), .A3(n119), .ZN(n79) );
  NAND2_X1 U18 ( .A1(A[6]), .A2(net56040), .ZN(n120) );
  NAND2_X1 U19 ( .A1(B[6]), .A2(net56046), .ZN(n121) );
  NAND2_X1 U20 ( .A1(F[6]), .A2(net56052), .ZN(n122) );
  AND3_X1 U21 ( .A1(n120), .A2(n121), .A3(n122), .ZN(n22) );
  NAND2_X1 U22 ( .A1(A[1]), .A2(net56036), .ZN(n123) );
  NAND2_X1 U23 ( .A1(B[1]), .A2(net56042), .ZN(n124) );
  NAND2_X1 U24 ( .A1(F[1]), .A2(net56048), .ZN(n125) );
  AND3_X1 U25 ( .A1(n123), .A2(n124), .A3(n125), .ZN(n73) );
  AND2_X1 U26 ( .A1(n133), .A2(n126), .ZN(n97) );
  NAND2_X1 U27 ( .A1(n19), .A2(n112), .ZN(Y[7]) );
  NAND2_X1 U28 ( .A1(n97), .A2(n110), .ZN(Y[12]) );
  NAND2_X1 U29 ( .A1(A[4]), .A2(net56040), .ZN(n127) );
  NAND2_X1 U30 ( .A1(B[4]), .A2(net56046), .ZN(n128) );
  NAND2_X1 U31 ( .A1(F[4]), .A2(net56052), .ZN(n129) );
  AND3_X1 U32 ( .A1(n127), .A2(n128), .A3(n129), .ZN(n28) );
  BUF_X1 U33 ( .A(n9), .Z(net56052) );
  AND2_X1 U34 ( .A1(n134), .A2(n135), .ZN(n130) );
  AND2_X1 U35 ( .A1(n136), .A2(n130), .ZN(n100) );
  NAND2_X1 U36 ( .A1(n100), .A2(n111), .ZN(Y[11]) );
  NAND2_X1 U37 ( .A1(A[12]), .A2(net56036), .ZN(n131) );
  NAND2_X1 U38 ( .A1(B[12]), .A2(net56042), .ZN(n132) );
  NAND2_X1 U39 ( .A1(F[12]), .A2(net56048), .ZN(n133) );
  NAND2_X1 U40 ( .A1(A[11]), .A2(net56036), .ZN(n134) );
  NAND2_X1 U41 ( .A1(B[11]), .A2(net56042), .ZN(n135) );
  NAND2_X1 U42 ( .A1(F[11]), .A2(net56048), .ZN(n136) );
  NAND2_X1 U43 ( .A1(A[7]), .A2(net56040), .ZN(n137) );
  NAND2_X1 U44 ( .A1(B[7]), .A2(net56046), .ZN(n138) );
  NAND2_X1 U45 ( .A1(F[7]), .A2(net56052), .ZN(n139) );
  AND3_X1 U46 ( .A1(n137), .A2(n138), .A3(n139), .ZN(n19) );
  NAND2_X1 U47 ( .A1(A[0]), .A2(net56036), .ZN(n140) );
  NAND2_X1 U48 ( .A1(B[0]), .A2(net56042), .ZN(n141) );
  NAND2_X1 U49 ( .A1(F[0]), .A2(net56048), .ZN(n142) );
  NAND2_X1 U50 ( .A1(n25), .A2(n113), .ZN(Y[5]) );
  NAND2_X1 U51 ( .A1(A[9]), .A2(net56040), .ZN(n143) );
  NAND2_X1 U52 ( .A1(B[9]), .A2(net56046), .ZN(n144) );
  NAND2_X1 U53 ( .A1(F[9]), .A2(net56052), .ZN(n145) );
  AND3_X1 U54 ( .A1(n143), .A2(n144), .A3(n145), .ZN(n6) );
  NAND2_X1 U55 ( .A1(A[2]), .A2(net56038), .ZN(n146) );
  NAND2_X1 U56 ( .A1(B[2]), .A2(net56044), .ZN(n147) );
  NAND2_X1 U57 ( .A1(F[2]), .A2(net56050), .ZN(n148) );
  AND3_X1 U58 ( .A1(n148), .A2(n147), .A3(n146), .ZN(n40) );
  AOI22_X1 U59 ( .A1(D[0]), .A2(net56054), .B1(H[0]), .B2(net56060), .ZN(n105)
         );
  NAND2_X1 U60 ( .A1(n105), .A2(n114), .ZN(Y[0]) );
  BUF_X1 U61 ( .A(n11), .Z(net56060) );
  BUF_X1 U62 ( .A(n10), .Z(net56054) );
  AND3_X1 U63 ( .A1(sel[1]), .A2(sel[0]), .A3(n107), .ZN(n11) );
  BUF_X1 U64 ( .A(n11), .Z(net56062) );
  BUF_X1 U65 ( .A(n11), .Z(net56064) );
  AND3_X1 U66 ( .A1(sel[0]), .A2(n108), .A3(sel[1]), .ZN(n10) );
  BUF_X1 U67 ( .A(n10), .Z(net56056) );
  BUF_X1 U68 ( .A(n10), .Z(net56058) );
  AND3_X1 U69 ( .A1(n108), .A2(net52587), .A3(sel[1]), .ZN(n13) );
  INV_X1 U70 ( .A(sel[1]), .ZN(n149) );
  AND3_X1 U71 ( .A1(net52587), .A2(n149), .A3(n107), .ZN(n12) );
  AND3_X1 U72 ( .A1(sel[0]), .A2(n149), .A3(n107), .ZN(n9) );
  AND3_X1 U73 ( .A1(net52587), .A2(n149), .A3(n108), .ZN(n7) );
  AND3_X1 U74 ( .A1(n108), .A2(n149), .A3(sel[0]), .ZN(n8) );
  NAND2_X1 U75 ( .A1(n32), .A2(n109), .ZN(Y[31]) );
  NAND2_X1 U76 ( .A1(A[5]), .A2(net56040), .ZN(n150) );
  NAND2_X1 U77 ( .A1(B[5]), .A2(net56046), .ZN(n151) );
  NAND2_X1 U78 ( .A1(F[5]), .A2(net56052), .ZN(n152) );
  AND3_X1 U79 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n25) );
  BUF_X1 U80 ( .A(n12), .Z(net56066) );
  BUF_X1 U81 ( .A(n12), .Z(net56068) );
  BUF_X1 U82 ( .A(n7), .Z(net56038) );
  BUF_X1 U83 ( .A(n7), .Z(net56036) );
  BUF_X1 U84 ( .A(n12), .Z(net56070) );
  BUF_X1 U85 ( .A(n7), .Z(net56040) );
  BUF_X1 U86 ( .A(n13), .Z(net56072) );
  BUF_X1 U87 ( .A(n13), .Z(net56074) );
  BUF_X1 U88 ( .A(n8), .Z(net56044) );
  BUF_X1 U89 ( .A(n8), .Z(net56042) );
  BUF_X1 U90 ( .A(n13), .Z(net56076) );
  BUF_X1 U91 ( .A(n8), .Z(net56046) );
  AOI222_X1 U92 ( .A1(A[3]), .A2(net56040), .B1(B[3]), .B2(net56046), .C1(F[3]), .C2(net56052), .ZN(n31) );
  AOI222_X1 U93 ( .A1(A[8]), .A2(net56040), .B1(B[8]), .B2(net56046), .C1(F[8]), .C2(net56052), .ZN(n16) );
  AOI222_X1 U94 ( .A1(A[31]), .A2(net56040), .B1(B[31]), .B2(net56046), .C1(
        F[31]), .C2(net56052), .ZN(n34) );
  AOI222_X1 U95 ( .A1(A[17]), .A2(net56036), .B1(B[17]), .B2(net56042), .C1(
        F[17]), .C2(net56048), .ZN(n82) );
  AOI222_X1 U96 ( .A1(A[14]), .A2(net56036), .B1(B[14]), .B2(net56042), .C1(
        F[14]), .C2(net56048), .ZN(n91) );
  AOI222_X1 U97 ( .A1(A[28]), .A2(net56038), .B1(B[28]), .B2(net56044), .C1(
        F[28]), .C2(net56050), .ZN(n46) );
  AOI222_X1 U98 ( .A1(A[23]), .A2(net56038), .B1(B[23]), .B2(net56044), .C1(
        F[23]), .C2(net56050), .ZN(n61) );
  AOI222_X1 U99 ( .A1(A[15]), .A2(net56036), .B1(B[15]), .B2(net56042), .C1(
        F[15]), .C2(net56048), .ZN(n88) );
  AOI222_X1 U100 ( .A1(A[27]), .A2(net56038), .B1(B[27]), .B2(net56044), .C1(
        F[27]), .C2(net56050), .ZN(n49) );
  AOI222_X1 U101 ( .A1(A[16]), .A2(net56036), .B1(B[16]), .B2(net56042), .C1(
        F[16]), .C2(net56048), .ZN(n85) );
  AOI222_X1 U102 ( .A1(A[24]), .A2(net56038), .B1(B[24]), .B2(net56044), .C1(
        F[24]), .C2(net56050), .ZN(n58) );
  AOI222_X1 U103 ( .A1(A[21]), .A2(net56038), .B1(B[21]), .B2(net56044), .C1(
        F[21]), .C2(net56050), .ZN(n67) );
  AOI222_X1 U104 ( .A1(A[10]), .A2(net56036), .B1(B[10]), .B2(net56042), .C1(
        F[10]), .C2(net56048), .ZN(n103) );
  AOI222_X1 U105 ( .A1(A[25]), .A2(net56038), .B1(B[25]), .B2(net56044), .C1(
        F[25]), .C2(net56050), .ZN(n55) );
  AOI222_X1 U106 ( .A1(A[22]), .A2(net56038), .B1(B[22]), .B2(net56044), .C1(
        F[22]), .C2(net56050), .ZN(n64) );
  AOI222_X1 U107 ( .A1(A[19]), .A2(net56036), .B1(B[19]), .B2(net56042), .C1(
        F[19]), .C2(net56048), .ZN(n76) );
  AOI222_X1 U108 ( .A1(A[20]), .A2(net56038), .B1(B[20]), .B2(net56044), .C1(
        F[20]), .C2(net56050), .ZN(n70) );
  AOI222_X1 U109 ( .A1(A[13]), .A2(net56036), .B1(B[13]), .B2(net56042), .C1(
        F[13]), .C2(net56048), .ZN(n94) );
  AOI222_X1 U112 ( .A1(A[26]), .A2(net56038), .B1(B[26]), .B2(net56044), .C1(
        F[26]), .C2(net56050), .ZN(n52) );
  AOI222_X1 U114 ( .A1(A[29]), .A2(net56038), .B1(B[29]), .B2(net56044), .C1(
        F[29]), .C2(net56050), .ZN(n43) );
  AOI222_X1 U117 ( .A1(A[30]), .A2(net56038), .B1(B[30]), .B2(net56044), .C1(
        F[30]), .C2(net56050), .ZN(n37) );
  AOI22_X1 U138 ( .A1(D[5]), .A2(net56058), .B1(H[5]), .B2(net56064), .ZN(n24)
         );
  AOI22_X1 U139 ( .A1(E[0]), .A2(net56066), .B1(C[0]), .B2(net56072), .ZN(n104) );
  AOI22_X1 U141 ( .A1(D[31]), .A2(net56058), .B1(H[31]), .B2(net56064), .ZN(
        n33) );
  AOI22_X1 U142 ( .A1(D[12]), .A2(net56054), .B1(H[12]), .B2(net56060), .ZN(
        n96) );
  AOI22_X1 U143 ( .A1(D[28]), .A2(net56056), .B1(H[28]), .B2(net56062), .ZN(
        n45) );
  AOI22_X1 U144 ( .A1(D[30]), .A2(net56056), .B1(H[30]), .B2(net56062), .ZN(
        n36) );
  AOI22_X1 U145 ( .A1(D[7]), .A2(net56058), .B1(H[7]), .B2(net56064), .ZN(n18)
         );
  AOI22_X1 U146 ( .A1(D[17]), .A2(net56054), .B1(H[17]), .B2(net56060), .ZN(
        n81) );
  AOI22_X1 U147 ( .A1(D[2]), .A2(net56056), .B1(H[2]), .B2(net56062), .ZN(n39)
         );
  AOI22_X1 U148 ( .A1(D[21]), .A2(net56056), .B1(H[21]), .B2(net56062), .ZN(
        n66) );
  AOI22_X1 U149 ( .A1(D[9]), .A2(net56058), .B1(H[9]), .B2(net56064), .ZN(n5)
         );
  AOI22_X1 U150 ( .A1(D[14]), .A2(net56054), .B1(H[14]), .B2(net56060), .ZN(
        n90) );
  AOI22_X1 U151 ( .A1(D[6]), .A2(net56058), .B1(H[6]), .B2(net56064), .ZN(n21)
         );
  AOI22_X1 U152 ( .A1(D[20]), .A2(net56056), .B1(H[20]), .B2(net56062), .ZN(
        n69) );
  AOI22_X1 U153 ( .A1(D[4]), .A2(net56058), .B1(H[4]), .B2(net56064), .ZN(n27)
         );
  AOI22_X1 U154 ( .A1(D[23]), .A2(net56056), .B1(H[23]), .B2(net56062), .ZN(
        n60) );
  AOI22_X1 U155 ( .A1(D[11]), .A2(net56054), .B1(H[11]), .B2(net56060), .ZN(
        n99) );
  AOI22_X1 U156 ( .A1(D[18]), .A2(net56054), .B1(H[18]), .B2(net56060), .ZN(
        n78) );
  AOI22_X1 U157 ( .A1(D[29]), .A2(net56056), .B1(H[29]), .B2(net56062), .ZN(
        n42) );
  AOI22_X1 U158 ( .A1(D[1]), .A2(net56054), .B1(H[1]), .B2(net56060), .ZN(n72)
         );
  AOI22_X1 U159 ( .A1(D[15]), .A2(net56054), .B1(H[15]), .B2(net56060), .ZN(
        n87) );
  AOI22_X1 U160 ( .A1(D[25]), .A2(net56056), .B1(H[25]), .B2(net56062), .ZN(
        n54) );
  AOI22_X1 U161 ( .A1(D[27]), .A2(net56056), .B1(H[27]), .B2(net56062), .ZN(
        n48) );
  AOI22_X1 U162 ( .A1(D[26]), .A2(net56056), .B1(H[26]), .B2(net56062), .ZN(
        n51) );
  AOI22_X1 U163 ( .A1(D[16]), .A2(net56054), .B1(H[16]), .B2(net56060), .ZN(
        n84) );
  AOI22_X1 U164 ( .A1(D[24]), .A2(net56056), .B1(H[24]), .B2(net56062), .ZN(
        n57) );
  AOI22_X1 U165 ( .A1(D[10]), .A2(net56054), .B1(H[10]), .B2(net56060), .ZN(
        n102) );
  AOI22_X1 U166 ( .A1(D[3]), .A2(net56058), .B1(H[3]), .B2(net56064), .ZN(n30)
         );
  AOI22_X1 U167 ( .A1(D[22]), .A2(net56056), .B1(H[22]), .B2(net56062), .ZN(
        n63) );
  AOI22_X1 U168 ( .A1(D[19]), .A2(net56054), .B1(H[19]), .B2(net56060), .ZN(
        n75) );
  AOI22_X1 U169 ( .A1(D[8]), .A2(net56058), .B1(H[8]), .B2(net56064), .ZN(n15)
         );
  AOI22_X1 U170 ( .A1(D[13]), .A2(net56054), .B1(H[13]), .B2(net56060), .ZN(
        n93) );
  AOI22_X1 U171 ( .A1(E[6]), .A2(net56070), .B1(C[6]), .B2(net56076), .ZN(n20)
         );
  AOI22_X1 U172 ( .A1(E[7]), .A2(net56070), .B1(C[7]), .B2(net56076), .ZN(n17)
         );
  AOI22_X1 U173 ( .A1(E[9]), .A2(net56070), .B1(C[9]), .B2(net56076), .ZN(n4)
         );
  AOI22_X1 U174 ( .A1(E[8]), .A2(net56070), .B1(C[8]), .B2(net56076), .ZN(n14)
         );
  AOI22_X1 U175 ( .A1(E[5]), .A2(net56070), .B1(C[5]), .B2(net56076), .ZN(n23)
         );
  AOI22_X1 U176 ( .A1(E[3]), .A2(net56070), .B1(C[3]), .B2(net56076), .ZN(n29)
         );
  AOI22_X1 U177 ( .A1(E[30]), .A2(net56068), .B1(C[30]), .B2(net56074), .ZN(
        n35) );
  AOI22_X1 U178 ( .A1(E[21]), .A2(net56068), .B1(C[21]), .B2(net56074), .ZN(
        n65) );
  AOI22_X1 U179 ( .A1(E[28]), .A2(net56068), .B1(C[28]), .B2(net56074), .ZN(
        n44) );
  AOI22_X1 U180 ( .A1(E[20]), .A2(net56068), .B1(C[20]), .B2(net56074), .ZN(
        n68) );
  AOI22_X1 U181 ( .A1(E[29]), .A2(net56068), .B1(C[29]), .B2(net56074), .ZN(
        n41) );
  AOI22_X1 U182 ( .A1(E[25]), .A2(net56068), .B1(C[25]), .B2(net56074), .ZN(
        n53) );
  AOI22_X1 U183 ( .A1(E[26]), .A2(net56068), .B1(C[26]), .B2(net56074), .ZN(
        n50) );
  AOI22_X1 U184 ( .A1(E[27]), .A2(net56068), .B1(C[27]), .B2(net56074), .ZN(
        n47) );
  AOI22_X1 U185 ( .A1(E[22]), .A2(net56068), .B1(C[22]), .B2(net56074), .ZN(
        n62) );
  AOI22_X1 U186 ( .A1(E[2]), .A2(net56068), .B1(C[2]), .B2(net56074), .ZN(n38)
         );
  AOI22_X1 U187 ( .A1(E[23]), .A2(net56068), .B1(C[23]), .B2(net56074), .ZN(
        n59) );
  AOI22_X1 U188 ( .A1(E[24]), .A2(net56068), .B1(C[24]), .B2(net56074), .ZN(
        n56) );
  AOI22_X1 U189 ( .A1(E[15]), .A2(net56066), .B1(C[15]), .B2(net56072), .ZN(
        n86) );
  AOI22_X1 U190 ( .A1(E[10]), .A2(net56066), .B1(C[10]), .B2(net56072), .ZN(
        n101) );
  AOI22_X1 U191 ( .A1(E[13]), .A2(net56066), .B1(C[13]), .B2(net56072), .ZN(
        n92) );
  AOI22_X1 U192 ( .A1(E[14]), .A2(net56066), .B1(C[14]), .B2(net56072), .ZN(
        n89) );
  AOI22_X1 U193 ( .A1(E[11]), .A2(net56066), .B1(C[11]), .B2(net56072), .ZN(
        n98) );
  AOI22_X1 U194 ( .A1(E[16]), .A2(net56066), .B1(C[16]), .B2(net56072), .ZN(
        n83) );
  AOI22_X1 U195 ( .A1(E[12]), .A2(net56066), .B1(C[12]), .B2(net56072), .ZN(
        n95) );
  AOI22_X1 U196 ( .A1(E[17]), .A2(net56066), .B1(C[17]), .B2(net56072), .ZN(
        n80) );
  AOI22_X1 U197 ( .A1(E[18]), .A2(net56066), .B1(C[18]), .B2(net56072), .ZN(
        n77) );
  AOI22_X1 U198 ( .A1(E[19]), .A2(net56066), .B1(C[19]), .B2(net56072), .ZN(
        n74) );
  AOI22_X1 U199 ( .A1(E[1]), .A2(net56066), .B1(C[1]), .B2(net56072), .ZN(n71)
         );
  NOR2_X1 U200 ( .A1(sel[2]), .A2(sel[3]), .ZN(n108) );
  NOR2_X1 U201 ( .A1(n153), .A2(sel[3]), .ZN(n107) );
  INV_X1 U202 ( .A(sel[2]), .ZN(n153) );
  INV_X1 U203 ( .A(sel[0]), .ZN(net52587) );
  AOI22_X1 U204 ( .A1(E[31]), .A2(net56070), .B1(C[31]), .B2(net56076), .ZN(
        n32) );
endmodule


module alu ( data_in1, data_in2, op_sel, data_out );
  input [31:0] data_in1;
  input [31:0] data_in2;
  input [3:0] op_sel;
  output [31:0] data_out;
  wire   p4_cin, add_sel, log_shift, N41, N42, N43, N44, N49, n54, n55, n56,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;
  wire   [3:0] mux_sel;
  wire   [2:0] cmp_sel;
  wire   [31:0] p4_operand;
  wire   [31:0] p4_out;
  wire   [31:0] and_out;
  wire   [31:0] or_out;
  wire   [31:0] xor_out;
  wire   [31:0] sl_out;
  wire   [31:0] sr_out;
  wire   [31:0] cmp_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  DLH_X1 \cmp_sel_reg[2]  ( .G(n121), .D(N49), .Q(cmp_sel[2]) );
  DLH_X1 \cmp_sel_reg[1]  ( .G(n121), .D(n55), .Q(cmp_sel[1]) );
  DLH_X1 \cmp_sel_reg[0]  ( .G(n121), .D(n54), .Q(cmp_sel[0]) );
  DLH_X1 p4_cin_reg ( .G(N41), .D(n56), .Q(p4_cin) );
  DLH_X1 \mux_sel_reg[2]  ( .G(N42), .D(n50), .Q(mux_sel[2]) );
  DLH_X1 \mux_sel_reg[1]  ( .G(N42), .D(N44), .Q(mux_sel[1]) );
  DLH_X1 \mux_sel_reg[0]  ( .G(N42), .D(N43), .Q(mux_sel[0]) );
  DLH_X1 log_shift_reg ( .G(n123), .D(n51), .Q(log_shift) );
  NAND3_X1 U57 ( .A1(n42), .A2(n40), .A3(n43), .ZN(N44) );
  NAND3_X1 U58 ( .A1(n42), .A2(n122), .A3(n44), .ZN(N42) );
  XOR2_X1 U59 ( .A(op_sel[2]), .B(op_sel[0]), .Z(n46) );
  XOR2_X1 U60 ( .A(op_sel[1]), .B(op_sel[0]), .Z(n49) );
  NAND3_X1 U61 ( .A1(n127), .A2(n126), .A3(op_sel[2]), .ZN(n42) );
  MUX21_GENERIC_NBIT32_2 mux_p4 ( .A({data_in2[31], n61, n78, n64, 
        data_in2[27], n62, data_in2[25], n52, n60, n57, n75, data_in2[20], n73, 
        data_in2[18:14], n53, data_in2[12:11], n58, n77, n76, n59, n74, 
        data_in2[5:4], n63, n70, n68, n72}), .B({n89, n90, n91, n92, n93, n94, 
        n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
        n119, n120}), .SEL(add_sel), .Y(p4_operand) );
  P4_ADDER_NBIT32_NBIT_PER_BLOCK4_1 add ( .A({data_in1[31], n88, 
        data_in1[29:23], n87, n86, data_in1[20:19], n85, data_in1[17:15], n84, 
        n83, data_in1[12:10], n82, n81, data_in1[7:5], n80, data_in1[3], n67, 
        n66, n79}), .B(p4_operand), .Cin(p4_cin), .Y(p4_out) );
  and_gate_nbit32 and_m ( .A({data_in1[31], n88, data_in1[29:23], n87, n86, 
        data_in1[20:19], n85, data_in1[17:15], n84, n83, data_in1[12:10], n82, 
        n81, data_in1[7:5], n80, data_in1[3], n67, n66, n79}), .B({
        data_in2[31], n61, n78, n64, data_in2[27], n62, data_in2[25], n52, n60, 
        n57, n75, data_in2[20], n73, data_in2[18:14], n53, data_in2[12:11], 
        n58, n77, n76, n59, n74, data_in2[5:4], n63, n71, n69, n72}), .Y(
        and_out) );
  or_gate_nbit32 or_m ( .A({data_in1[31], n88, data_in1[29:23], n87, n86, 
        data_in1[20:19], n85, data_in1[17:15], n84, n83, data_in1[12:10], n82, 
        n81, data_in1[7:5], n80, data_in1[3], n67, n66, n79}), .B({
        data_in2[31], n61, n78, n64, data_in2[27], n62, data_in2[25], n52, n60, 
        n57, n75, data_in2[20], n73, data_in2[18:14], n53, data_in2[12:11], 
        n58, n77, n76, n59, n74, data_in2[5:4], n63, n71, n69, n72}), .Y(
        or_out) );
  xor_gate_nbit32 xor_m ( .A({data_in1[31], n88, data_in1[29:23], n87, n86, 
        data_in1[20:19], n85, data_in1[17:15], n84, n83, data_in1[12:10], n82, 
        n81, data_in1[7:5], n80, data_in1[3], n67, n66, n79}), .B({
        data_in2[31], n61, n78, n64, data_in2[27], n62, data_in2[25], n52, n60, 
        n57, n75, data_in2[20], n73, data_in2[18:14], n53, data_in2[12:11], 
        n58, n77, n76, n59, n74, data_in2[5:4], n63, n70, n68, n72}), .Y(
        xor_out) );
  shifter_sx_nbit32 sl ( .r1({data_in1[31], n88, data_in1[29:23], n87, n86, 
        data_in1[20:19], n85, data_in1[17:15], n84, n83, data_in1[12:10], n82, 
        n81, data_in1[7:5], n80, data_in1[3], n67, n66, n79}), .r2({
        data_in2[31:4], n63, n71, n69, n72}), .data_out(sl_out) );
  shifter_dx_nbit32 sr ( .r1({data_in1[31], n88, data_in1[29:23], n87, n86, 
        data_in1[20:19], n85, data_in1[17:15], n84, n83, data_in1[12:10], n82, 
        n81, data_in1[7:5], n80, data_in1[3], n67, n66, n79}), .r2({
        data_in2[31], n61, data_in2[29:11], n58, data_in2[9:4], n63, n70, n68, 
        n72}), .log(log_shift), .data_out(sr_out) );
  comparator cmp ( .r1({data_in1[31], n88, data_in1[29:23], n87, n86, 
        data_in1[20:19], n85, data_in1[17:15], n84, n83, data_in1[12:10], n82, 
        n81, data_in1[7:5], n80, data_in1[3:0]}), .r2({data_in2[31], n61, n78, 
        n64, data_in2[27], n62, data_in2[25], n52, n60, n57, n75, data_in2[20], 
        n73, data_in2[18:14], n53, data_in2[12:11], n58, n77, n76, n59, n74, 
        data_in2[5:0]}), .sel(cmp_sel), .data_out({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, cmp_out[0]}) );
  mux11to1_nbit32 mux ( .A(p4_out), .B(and_out), .C(or_out), .D(xor_out), .E(
        sl_out), .F(sr_out), .H({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        cmp_out[0]}), .sel({1'b0, mux_sel[2:0]}), .Y(data_out) );
  DLH_X1 add_sel_reg ( .G(N41), .D(n56), .Q(add_sel) );
  BUF_X1 U3 ( .A(n65), .Z(n71) );
  BUF_X2 U4 ( .A(data_in2[3]), .Z(n63) );
  BUF_X1 U5 ( .A(data_in1[13]), .Z(n83) );
  BUF_X1 U6 ( .A(data_in1[14]), .Z(n84) );
  BUF_X2 U7 ( .A(data_in1[18]), .Z(n85) );
  NOR4_X1 U8 ( .A1(n45), .A2(N49), .A3(n54), .A4(n55), .ZN(n40) );
  BUF_X1 U9 ( .A(data_in1[9]), .Z(n82) );
  CLKBUF_X1 U10 ( .A(data_in2[24]), .Z(n52) );
  CLKBUF_X1 U11 ( .A(data_in2[13]), .Z(n53) );
  CLKBUF_X1 U12 ( .A(data_in2[22]), .Z(n57) );
  BUF_X2 U13 ( .A(data_in2[10]), .Z(n58) );
  CLKBUF_X1 U14 ( .A(data_in2[7]), .Z(n59) );
  CLKBUF_X1 U15 ( .A(data_in2[23]), .Z(n60) );
  BUF_X1 U16 ( .A(data_in2[2]), .Z(n65) );
  BUF_X2 U17 ( .A(data_in2[30]), .Z(n61) );
  CLKBUF_X1 U18 ( .A(data_in2[26]), .Z(n62) );
  CLKBUF_X1 U19 ( .A(data_in2[28]), .Z(n64) );
  CLKBUF_X1 U20 ( .A(data_in1[1]), .Z(n66) );
  CLKBUF_X1 U21 ( .A(data_in1[0]), .Z(n79) );
  CLKBUF_X1 U22 ( .A(data_in2[0]), .Z(n72) );
  INV_X1 U23 ( .A(n69), .ZN(n119) );
  INV_X1 U24 ( .A(n77), .ZN(n111) );
  INV_X1 U25 ( .A(n74), .ZN(n114) );
  INV_X1 U26 ( .A(n71), .ZN(n118) );
  INV_X1 U27 ( .A(n73), .ZN(n101) );
  INV_X1 U28 ( .A(n78), .ZN(n91) );
  INV_X1 U29 ( .A(n58), .ZN(n110) );
  INV_X1 U30 ( .A(n63), .ZN(n117) );
  INV_X1 U31 ( .A(n62), .ZN(n94) );
  INV_X1 U32 ( .A(data_in2[4]), .ZN(n116) );
  INV_X1 U33 ( .A(data_in2[31]), .ZN(n89) );
  INV_X1 U34 ( .A(data_in2[11]), .ZN(n109) );
  INV_X1 U35 ( .A(data_in2[12]), .ZN(n108) );
  INV_X1 U36 ( .A(data_in2[14]), .ZN(n106) );
  INV_X1 U37 ( .A(data_in2[15]), .ZN(n105) );
  INV_X1 U38 ( .A(n60), .ZN(n97) );
  INV_X1 U39 ( .A(data_in2[17]), .ZN(n103) );
  INV_X1 U40 ( .A(data_in2[16]), .ZN(n104) );
  INV_X1 U41 ( .A(data_in2[18]), .ZN(n102) );
  INV_X1 U42 ( .A(data_in2[5]), .ZN(n115) );
  INV_X1 U43 ( .A(n61), .ZN(n90) );
  INV_X1 U44 ( .A(data_in2[27]), .ZN(n93) );
  INV_X1 U45 ( .A(data_in2[25]), .ZN(n95) );
  INV_X1 U46 ( .A(data_in2[20]), .ZN(n100) );
  INV_X1 U47 ( .A(n59), .ZN(n113) );
  INV_X1 U48 ( .A(n52), .ZN(n96) );
  NOR2_X1 U49 ( .A1(n124), .A2(n42), .ZN(n55) );
  OR3_X1 U50 ( .A1(n126), .A2(n127), .A3(n44), .ZN(n43) );
  INV_X1 U51 ( .A(n40), .ZN(n121) );
  INV_X1 U52 ( .A(n50), .ZN(n122) );
  NAND2_X1 U53 ( .A1(n41), .A2(n40), .ZN(n50) );
  NAND2_X1 U54 ( .A1(n125), .A2(n124), .ZN(n44) );
  INV_X1 U55 ( .A(n41), .ZN(n123) );
  BUF_X1 U56 ( .A(data_in1[21]), .Z(n86) );
  BUF_X1 U93 ( .A(data_in1[22]), .Z(n87) );
  BUF_X1 U94 ( .A(data_in1[30]), .Z(n88) );
  AND2_X1 U95 ( .A1(n47), .A2(op_sel[1]), .ZN(n45) );
  NOR4_X1 U96 ( .A1(n127), .A2(n124), .A3(n125), .A4(op_sel[1]), .ZN(n54) );
  AOI211_X1 U97 ( .C1(n126), .C2(n47), .A(n48), .B(n51), .ZN(n41) );
  NOR3_X1 U98 ( .A1(n125), .A2(op_sel[3]), .A3(n127), .ZN(n48) );
  NOR3_X1 U99 ( .A1(op_sel[0]), .A2(op_sel[2]), .A3(n124), .ZN(n47) );
  NOR2_X1 U100 ( .A1(n44), .A2(op_sel[1]), .ZN(N41) );
  INV_X1 U101 ( .A(op_sel[3]), .ZN(n124) );
  INV_X1 U102 ( .A(op_sel[0]), .ZN(n127) );
  INV_X1 U103 ( .A(op_sel[2]), .ZN(n125) );
  INV_X1 U104 ( .A(op_sel[1]), .ZN(n126) );
  OAI21_X1 U105 ( .B1(op_sel[0]), .B2(N41), .A(n40), .ZN(N43) );
  AND3_X1 U106 ( .A1(op_sel[3]), .A2(n46), .A3(op_sel[1]), .ZN(N49) );
  AND3_X1 U107 ( .A1(n49), .A2(n124), .A3(op_sel[2]), .ZN(n51) );
  AND2_X1 U108 ( .A1(op_sel[0]), .A2(N41), .ZN(n56) );
  CLKBUF_X1 U109 ( .A(data_in1[2]), .Z(n67) );
  INV_X1 U110 ( .A(n53), .ZN(n107) );
  CLKBUF_X1 U111 ( .A(data_in2[1]), .Z(n68) );
  CLKBUF_X1 U112 ( .A(data_in2[1]), .Z(n69) );
  CLKBUF_X1 U113 ( .A(n65), .Z(n70) );
  CLKBUF_X1 U114 ( .A(data_in2[19]), .Z(n73) );
  CLKBUF_X1 U115 ( .A(data_in2[6]), .Z(n74) );
  CLKBUF_X1 U116 ( .A(data_in2[21]), .Z(n75) );
  INV_X1 U117 ( .A(n57), .ZN(n98) );
  CLKBUF_X1 U118 ( .A(data_in2[8]), .Z(n76) );
  CLKBUF_X1 U119 ( .A(data_in2[9]), .Z(n77) );
  CLKBUF_X1 U120 ( .A(data_in2[29]), .Z(n78) );
  INV_X1 U121 ( .A(n64), .ZN(n92) );
  INV_X1 U122 ( .A(n75), .ZN(n99) );
  INV_X1 U123 ( .A(n72), .ZN(n120) );
  INV_X1 U124 ( .A(n76), .ZN(n112) );
  CLKBUF_X3 U125 ( .A(data_in1[4]), .Z(n80) );
  CLKBUF_X3 U126 ( .A(data_in1[8]), .Z(n81) );
endmodule


module REG_GEN_NBIT32_9 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, net52311, net52312, net52338,
         net54370, net54368, net54366, net54364, net54362, net54360, net54356,
         net54354, net54352, net54350, net54498, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100,
         n101, n102, n103;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n41), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n43), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n43), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n43), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n43), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n42), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n43), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n42), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n42), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n42), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n42), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n43), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n42), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n42), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n43), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n42), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n42), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n42), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n41), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n42), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n41), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n41), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n41), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n41), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n41), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n41), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n41), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n41), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n41), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n41), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n42), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n43), .Q(Q[0]), .QN(n97) );
  OAI22_X1 U2 ( .A1(n97), .A2(net54354), .B1(n36), .B2(n37), .ZN(n35) );
  BUF_X1 U3 ( .A(n39), .Z(n37) );
  OAI22_X1 U4 ( .A1(n67), .A2(net54354), .B1(n37), .B2(net52311), .ZN(n5) );
  OAI22_X1 U5 ( .A1(n96), .A2(net54354), .B1(n37), .B2(net52338), .ZN(n34) );
  OAI22_X1 U6 ( .A1(n66), .A2(net54354), .B1(net52312), .B2(n37), .ZN(n4) );
  BUF_X1 U7 ( .A(Enable_n), .Z(n39) );
  BUF_X1 U8 ( .A(n39), .Z(net54356) );
  BUF_X1 U9 ( .A(n39), .Z(net54360) );
  INV_X1 U10 ( .A(D[0]), .ZN(n36) );
  INV_X1 U11 ( .A(n38), .ZN(net54354) );
  BUF_X1 U12 ( .A(n40), .Z(n38) );
  INV_X1 U13 ( .A(n38), .ZN(net54350) );
  INV_X1 U14 ( .A(n38), .ZN(net54352) );
  BUF_X1 U15 ( .A(Enable_n), .Z(n40) );
  BUF_X1 U16 ( .A(n40), .Z(net54368) );
  BUF_X1 U17 ( .A(n40), .Z(net54370) );
  BUF_X1 U18 ( .A(Enable_n), .Z(net54498) );
  BUF_X1 U19 ( .A(RESET_n), .Z(n42) );
  BUF_X1 U20 ( .A(RESET_n), .Z(n41) );
  BUF_X1 U21 ( .A(RESET_n), .Z(n43) );
  BUF_X1 U22 ( .A(net54498), .Z(net54362) );
  BUF_X1 U23 ( .A(net54498), .Z(net54366) );
  BUF_X1 U24 ( .A(net54498), .Z(net54364) );
  INV_X1 U25 ( .A(D[28]), .ZN(n103) );
  INV_X1 U26 ( .A(D[30]), .ZN(net52311) );
  OAI22_X1 U27 ( .A1(n90), .A2(net54352), .B1(net54362), .B2(n46), .ZN(n28) );
  INV_X1 U28 ( .A(D[7]), .ZN(n46) );
  OAI22_X1 U29 ( .A1(n80), .A2(net54350), .B1(net54366), .B2(n60), .ZN(n18) );
  INV_X1 U30 ( .A(D[17]), .ZN(n60) );
  OAI22_X1 U31 ( .A1(n95), .A2(net54352), .B1(n45), .B2(net54360), .ZN(n33) );
  INV_X1 U32 ( .A(D[2]), .ZN(n45) );
  OAI22_X1 U33 ( .A1(n76), .A2(net54350), .B1(net54368), .B2(n64), .ZN(n14) );
  INV_X1 U34 ( .A(D[21]), .ZN(n64) );
  OAI22_X1 U35 ( .A1(n88), .A2(net54352), .B1(net54362), .B2(n52), .ZN(n26) );
  INV_X1 U36 ( .A(D[9]), .ZN(n52) );
  OAI22_X1 U37 ( .A1(n83), .A2(net54350), .B1(n55), .B2(net54366), .ZN(n21) );
  INV_X1 U38 ( .A(D[14]), .ZN(n55) );
  OAI22_X1 U39 ( .A1(n91), .A2(net54352), .B1(n47), .B2(net54362), .ZN(n29) );
  INV_X1 U40 ( .A(D[6]), .ZN(n47) );
  OAI22_X1 U41 ( .A1(n77), .A2(net54350), .B1(net54368), .B2(n65), .ZN(n15) );
  INV_X1 U42 ( .A(D[20]), .ZN(n65) );
  OAI22_X1 U43 ( .A1(n93), .A2(net54352), .B1(net54360), .B2(n49), .ZN(n31) );
  INV_X1 U44 ( .A(D[4]), .ZN(n49) );
  OAI22_X1 U45 ( .A1(n74), .A2(net54350), .B1(net54370), .B2(n62), .ZN(n12) );
  INV_X1 U46 ( .A(D[23]), .ZN(n62) );
  OAI22_X1 U47 ( .A1(n86), .A2(net54352), .B1(net54364), .B2(n50), .ZN(n24) );
  INV_X1 U48 ( .A(D[11]), .ZN(n50) );
  OAI22_X1 U49 ( .A1(n79), .A2(net54350), .B1(n59), .B2(net54368), .ZN(n17) );
  INV_X1 U50 ( .A(D[18]), .ZN(n59) );
  OAI22_X1 U51 ( .A1(n68), .A2(net54354), .B1(net54356), .B2(n102), .ZN(n6) );
  INV_X1 U52 ( .A(D[29]), .ZN(n102) );
  INV_X1 U53 ( .A(D[1]), .ZN(net52338) );
  OAI22_X1 U54 ( .A1(n82), .A2(net54350), .B1(net54366), .B2(n54), .ZN(n20) );
  INV_X1 U55 ( .A(D[15]), .ZN(n54) );
  OAI22_X1 U56 ( .A1(n72), .A2(net54350), .B1(net54370), .B2(n100), .ZN(n10)
         );
  INV_X1 U57 ( .A(D[25]), .ZN(n100) );
  OAI22_X1 U58 ( .A1(n70), .A2(net54354), .B1(net54356), .B2(n98), .ZN(n8) );
  INV_X1 U59 ( .A(D[27]), .ZN(n98) );
  OAI22_X1 U60 ( .A1(n71), .A2(net54354), .B1(net54356), .B2(n99), .ZN(n9) );
  INV_X1 U61 ( .A(D[26]), .ZN(n99) );
  OAI22_X1 U62 ( .A1(n81), .A2(net54350), .B1(net54366), .B2(n61), .ZN(n19) );
  INV_X1 U63 ( .A(D[16]), .ZN(n61) );
  OAI22_X1 U64 ( .A1(n73), .A2(net54350), .B1(net54370), .B2(n101), .ZN(n11)
         );
  INV_X1 U65 ( .A(D[24]), .ZN(n101) );
  OAI22_X1 U66 ( .A1(n87), .A2(net54352), .B1(net54364), .B2(n51), .ZN(n25) );
  INV_X1 U67 ( .A(D[10]), .ZN(n51) );
  OAI22_X1 U68 ( .A1(n94), .A2(net54352), .B1(net54360), .B2(n44), .ZN(n32) );
  INV_X1 U69 ( .A(D[3]), .ZN(n44) );
  OAI22_X1 U70 ( .A1(n75), .A2(net54350), .B1(net54370), .B2(n63), .ZN(n13) );
  INV_X1 U71 ( .A(D[22]), .ZN(n63) );
  OAI22_X1 U72 ( .A1(n78), .A2(net54350), .B1(net54368), .B2(n58), .ZN(n16) );
  INV_X1 U73 ( .A(D[19]), .ZN(n58) );
  OAI22_X1 U74 ( .A1(n89), .A2(net54352), .B1(net54362), .B2(n53), .ZN(n27) );
  INV_X1 U75 ( .A(D[8]), .ZN(n53) );
  OAI22_X1 U76 ( .A1(n84), .A2(net54352), .B1(net54364), .B2(n56), .ZN(n22) );
  INV_X1 U77 ( .A(D[13]), .ZN(n56) );
  OAI22_X1 U78 ( .A1(n69), .A2(net54354), .B1(n103), .B2(net54356), .ZN(n7) );
  INV_X1 U79 ( .A(D[31]), .ZN(net52312) );
  OAI22_X1 U80 ( .A1(n85), .A2(net54352), .B1(n57), .B2(net54364), .ZN(n23) );
  INV_X1 U81 ( .A(D[12]), .ZN(n57) );
  INV_X1 U82 ( .A(D[5]), .ZN(n48) );
  OAI22_X1 U83 ( .A1(n92), .A2(net54352), .B1(n48), .B2(net54360), .ZN(n30) );
endmodule


module REG_GEN_NBIT32_8 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n52), .Q(Q[31]), .QN(n148) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n52), .Q(Q[30]), .QN(n147) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n52), .Q(Q[29]), .QN(n146) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n52), .Q(Q[28]), .QN(n145) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n52), .Q(Q[27]), .QN(n144) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n51), .Q(Q[26]), .QN(n143) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n51), .Q(Q[25]), .QN(n142) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n51), .Q(Q[24]), .QN(n141) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n51), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n51), .Q(Q[22]), .QN(n139) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n51), .Q(Q[21]), .QN(n138) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n52), .Q(Q[20]), .QN(n137) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n136) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n135) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n52), .Q(Q[17]), .QN(n134) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n133) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n132) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n131) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n50), .Q(Q[13]), .QN(n130) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n50), .Q(Q[12]), .QN(n129) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n50), .Q(Q[11]), .QN(n128) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n50), .Q(Q[10]), .QN(n127) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n50), .Q(Q[9]), .QN(n126) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n50), .Q(Q[8]), .QN(n125) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n50), .Q(Q[7]), .QN(n124) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n50), .Q(Q[6]), .QN(n123) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n50), .Q(Q[5]), .QN(n122) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n50), .Q(Q[4]), .QN(n121) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n50), .Q(Q[3]), .QN(n120) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n50), .Q(Q[2]), .QN(n119) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n51), .Q(Q[1]), .QN(n118) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n52), .Q(Q[0]), .QN(n117) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n44) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n146), .A2(n40), .B1(n41), .B2(n55), .ZN(n6) );
  INV_X1 U20 ( .A(D[29]), .ZN(n55) );
  OAI22_X1 U21 ( .A1(n117), .A2(n39), .B1(n42), .B2(n116), .ZN(n35) );
  INV_X1 U22 ( .A(D[0]), .ZN(n116) );
  OAI22_X1 U23 ( .A1(n118), .A2(n40), .B1(n42), .B2(n115), .ZN(n34) );
  INV_X1 U24 ( .A(D[1]), .ZN(n115) );
  OAI22_X1 U25 ( .A1(n143), .A2(n39), .B1(n41), .B2(n58), .ZN(n9) );
  INV_X1 U26 ( .A(D[26]), .ZN(n58) );
  OAI22_X1 U27 ( .A1(n144), .A2(n40), .B1(n41), .B2(n57), .ZN(n8) );
  INV_X1 U28 ( .A(D[27]), .ZN(n57) );
  OAI22_X1 U29 ( .A1(n145), .A2(n39), .B1(n41), .B2(n56), .ZN(n7) );
  OAI22_X1 U30 ( .A1(n147), .A2(n40), .B1(n42), .B2(n54), .ZN(n5) );
  INV_X1 U31 ( .A(D[30]), .ZN(n54) );
  OAI22_X1 U32 ( .A1(n148), .A2(n39), .B1(n42), .B2(n53), .ZN(n4) );
  INV_X1 U33 ( .A(D[31]), .ZN(n53) );
  OAI22_X1 U34 ( .A1(n119), .A2(n40), .B1(n43), .B2(n114), .ZN(n33) );
  INV_X1 U35 ( .A(D[2]), .ZN(n114) );
  OAI22_X1 U36 ( .A1(n120), .A2(n40), .B1(n43), .B2(n113), .ZN(n32) );
  INV_X1 U37 ( .A(D[3]), .ZN(n113) );
  OAI22_X1 U38 ( .A1(n121), .A2(n40), .B1(n43), .B2(n112), .ZN(n31) );
  INV_X1 U39 ( .A(D[4]), .ZN(n112) );
  OAI22_X1 U40 ( .A1(n122), .A2(n40), .B1(n43), .B2(n111), .ZN(n30) );
  INV_X1 U41 ( .A(D[5]), .ZN(n111) );
  OAI22_X1 U42 ( .A1(n123), .A2(n40), .B1(n44), .B2(n110), .ZN(n29) );
  INV_X1 U43 ( .A(D[6]), .ZN(n110) );
  OAI22_X1 U44 ( .A1(n124), .A2(n40), .B1(n44), .B2(n109), .ZN(n28) );
  INV_X1 U45 ( .A(D[7]), .ZN(n109) );
  OAI22_X1 U46 ( .A1(n125), .A2(n40), .B1(n44), .B2(n108), .ZN(n27) );
  INV_X1 U47 ( .A(D[8]), .ZN(n108) );
  OAI22_X1 U48 ( .A1(n126), .A2(n40), .B1(n44), .B2(n107), .ZN(n26) );
  INV_X1 U49 ( .A(D[9]), .ZN(n107) );
  OAI22_X1 U50 ( .A1(n127), .A2(n40), .B1(n45), .B2(n106), .ZN(n25) );
  INV_X1 U51 ( .A(D[10]), .ZN(n106) );
  OAI22_X1 U52 ( .A1(n128), .A2(n40), .B1(n45), .B2(n105), .ZN(n24) );
  INV_X1 U53 ( .A(D[11]), .ZN(n105) );
  OAI22_X1 U54 ( .A1(n129), .A2(n40), .B1(n45), .B2(n104), .ZN(n23) );
  INV_X1 U55 ( .A(D[12]), .ZN(n104) );
  OAI22_X1 U56 ( .A1(n130), .A2(n40), .B1(n45), .B2(n103), .ZN(n22) );
  INV_X1 U57 ( .A(D[13]), .ZN(n103) );
  OAI22_X1 U58 ( .A1(n131), .A2(n39), .B1(n46), .B2(n102), .ZN(n21) );
  INV_X1 U59 ( .A(D[14]), .ZN(n102) );
  OAI22_X1 U60 ( .A1(n132), .A2(n39), .B1(n46), .B2(n101), .ZN(n20) );
  INV_X1 U61 ( .A(D[15]), .ZN(n101) );
  OAI22_X1 U62 ( .A1(n133), .A2(n39), .B1(n46), .B2(n100), .ZN(n19) );
  INV_X1 U63 ( .A(D[16]), .ZN(n100) );
  OAI22_X1 U64 ( .A1(n134), .A2(n39), .B1(n46), .B2(n99), .ZN(n18) );
  INV_X1 U65 ( .A(D[17]), .ZN(n99) );
  OAI22_X1 U66 ( .A1(n135), .A2(n39), .B1(n47), .B2(n98), .ZN(n17) );
  INV_X1 U67 ( .A(D[18]), .ZN(n98) );
  OAI22_X1 U68 ( .A1(n136), .A2(n39), .B1(n47), .B2(n65), .ZN(n16) );
  OAI22_X1 U69 ( .A1(n137), .A2(n39), .B1(n47), .B2(n64), .ZN(n15) );
  INV_X1 U70 ( .A(D[20]), .ZN(n64) );
  OAI22_X1 U71 ( .A1(n138), .A2(n39), .B1(n47), .B2(n63), .ZN(n14) );
  INV_X1 U72 ( .A(D[21]), .ZN(n63) );
  OAI22_X1 U73 ( .A1(n139), .A2(n39), .B1(n48), .B2(n62), .ZN(n13) );
  OAI22_X1 U74 ( .A1(n140), .A2(n39), .B1(n48), .B2(n61), .ZN(n12) );
  INV_X1 U75 ( .A(D[23]), .ZN(n61) );
  OAI22_X1 U76 ( .A1(n141), .A2(n39), .B1(n48), .B2(n60), .ZN(n11) );
  INV_X1 U77 ( .A(D[24]), .ZN(n60) );
  OAI22_X1 U78 ( .A1(n142), .A2(n39), .B1(n48), .B2(n59), .ZN(n10) );
  INV_X1 U79 ( .A(D[25]), .ZN(n59) );
  INV_X1 U80 ( .A(D[28]), .ZN(n56) );
  INV_X1 U81 ( .A(D[19]), .ZN(n65) );
  INV_X1 U82 ( .A(D[22]), .ZN(n62) );
endmodule


module PG_block_96 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_30 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module PG_block_95 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_94 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_93 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_92 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_91 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_90 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_89 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_88 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_87 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_86 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_85 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_84 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_83 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_82 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_81 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_80 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_79 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_78 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_77 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_76 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_75 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_74 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_73 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_72 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_71 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_70 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_69 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_68 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_67 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_66 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_65 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_29 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_81 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_28 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_80 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_79 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_78 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_77 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_76 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_75 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_74 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_73 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_72 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_71 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_70 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_69 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_68 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_67 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_66 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_65 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_64 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_63 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_62 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_61 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_60 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_G_27 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_59 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_26 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_25 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_58 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_57 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_56 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_55 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_24 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_23 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_22 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_21 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   Cin, first_generate, \p_vett[4][3] , \p_vett[4][2] , \p_vett[3][3] ,
         \p_vett[3][2] , \p_vett[3][1] , \p_vett[2][7] , \p_vett[2][6] ,
         \p_vett[2][5] , \p_vett[2][4] , \p_vett[2][3] , \p_vett[2][2] ,
         \p_vett[2][1] , \p_vett[1][15] , \p_vett[1][14] , \p_vett[1][13] ,
         \p_vett[1][12] , \p_vett[1][11] , \p_vett[1][10] , \p_vett[1][9] ,
         \p_vett[1][8] , \p_vett[1][7] , \p_vett[1][6] , \p_vett[1][5] ,
         \p_vett[1][4] , \p_vett[1][3] , \p_vett[1][2] , \p_vett[1][1] ,
         \p_vett[0][31] , \p_vett[0][30] , \p_vett[0][29] , \p_vett[0][28] ,
         \p_vett[0][27] , \p_vett[0][26] , \p_vett[0][25] , \p_vett[0][24] ,
         \p_vett[0][23] , \p_vett[0][22] , \p_vett[0][21] , \p_vett[0][20] ,
         \p_vett[0][19] , \p_vett[0][18] , \p_vett[0][17] , \p_vett[0][16] ,
         \p_vett[0][15] , \p_vett[0][14] , \p_vett[0][13] , \p_vett[0][12] ,
         \p_vett[0][11] , \p_vett[0][10] , \p_vett[0][9] , \p_vett[0][8] ,
         \p_vett[0][7] , \p_vett[0][6] , \p_vett[0][5] , \p_vett[0][4] ,
         \p_vett[0][3] , \p_vett[0][2] , \p_vett[0][1] , \p_vett[0][0] ,
         \g_vett[4][3] , \g_vett[4][2] , \g_vett[3][3] , \g_vett[3][2] ,
         \g_vett[3][1] , \g_vett[2][7] , \g_vett[2][6] , \g_vett[2][5] ,
         \g_vett[2][4] , \g_vett[2][3] , \g_vett[2][2] , \g_vett[2][1] ,
         \g_vett[1][15] , \g_vett[1][14] , \g_vett[1][13] , \g_vett[1][12] ,
         \g_vett[1][11] , \g_vett[1][10] , \g_vett[1][9] , \g_vett[1][8] ,
         \g_vett[1][7] , \g_vett[1][6] , \g_vett[1][5] , \g_vett[1][4] ,
         \g_vett[1][3] , \g_vett[1][2] , \g_vett[1][1] , \g_vett[1][0] ,
         \g_vett[0][31] , \g_vett[0][30] , \g_vett[0][29] , \g_vett[0][28] ,
         \g_vett[0][27] , \g_vett[0][26] , \g_vett[0][25] , \g_vett[0][24] ,
         \g_vett[0][23] , \g_vett[0][22] , \g_vett[0][21] , \g_vett[0][20] ,
         \g_vett[0][19] , \g_vett[0][18] , \g_vett[0][17] , \g_vett[0][16] ,
         \g_vett[0][15] , \g_vett[0][14] , \g_vett[0][13] , \g_vett[0][12] ,
         \g_vett[0][11] , \g_vett[0][10] , \g_vett[0][9] , \g_vett[0][8] ,
         \g_vett[0][7] , \g_vett[0][6] , \g_vett[0][5] , \g_vett[0][4] ,
         \g_vett[0][3] , \g_vett[0][2] , \g_vett[0][1] , \g_vett[0][0] ;
  assign Co[0] = Cin;

  PG_block_96 PGblock_first ( .A(A[0]), .B(B[0]), .G(first_generate), .P(
        \p_vett[0][0] ) );
  GENERAL_G_30 G_first ( .G_in(first_generate), .P_in(\p_vett[0][0] ), 
        .G_in_prev(Cin), .G_out(\g_vett[0][0] ) );
  PG_block_95 PG_0_1 ( .A(A[1]), .B(B[1]), .G(\g_vett[0][1] ), .P(
        \p_vett[0][1] ) );
  PG_block_94 PG_0_2 ( .A(A[2]), .B(B[2]), .G(\g_vett[0][2] ), .P(
        \p_vett[0][2] ) );
  PG_block_93 PG_0_3 ( .A(A[3]), .B(B[3]), .G(\g_vett[0][3] ), .P(
        \p_vett[0][3] ) );
  PG_block_92 PG_0_4 ( .A(A[4]), .B(B[4]), .G(\g_vett[0][4] ), .P(
        \p_vett[0][4] ) );
  PG_block_91 PG_0_5 ( .A(A[5]), .B(B[5]), .G(\g_vett[0][5] ), .P(
        \p_vett[0][5] ) );
  PG_block_90 PG_0_6 ( .A(A[6]), .B(B[6]), .G(\g_vett[0][6] ), .P(
        \p_vett[0][6] ) );
  PG_block_89 PG_0_7 ( .A(A[7]), .B(B[7]), .G(\g_vett[0][7] ), .P(
        \p_vett[0][7] ) );
  PG_block_88 PG_0_8 ( .A(A[8]), .B(B[8]), .G(\g_vett[0][8] ), .P(
        \p_vett[0][8] ) );
  PG_block_87 PG_0_9 ( .A(A[9]), .B(B[9]), .G(\g_vett[0][9] ), .P(
        \p_vett[0][9] ) );
  PG_block_86 PG_0_10 ( .A(A[10]), .B(B[10]), .G(\g_vett[0][10] ), .P(
        \p_vett[0][10] ) );
  PG_block_85 PG_0_11 ( .A(A[11]), .B(B[11]), .G(\g_vett[0][11] ), .P(
        \p_vett[0][11] ) );
  PG_block_84 PG_0_12 ( .A(A[12]), .B(B[12]), .G(\g_vett[0][12] ), .P(
        \p_vett[0][12] ) );
  PG_block_83 PG_0_13 ( .A(A[13]), .B(B[13]), .G(\g_vett[0][13] ), .P(
        \p_vett[0][13] ) );
  PG_block_82 PG_0_14 ( .A(A[14]), .B(B[14]), .G(\g_vett[0][14] ), .P(
        \p_vett[0][14] ) );
  PG_block_81 PG_0_15 ( .A(A[15]), .B(B[15]), .G(\g_vett[0][15] ), .P(
        \p_vett[0][15] ) );
  PG_block_80 PG_0_16 ( .A(A[16]), .B(B[16]), .G(\g_vett[0][16] ), .P(
        \p_vett[0][16] ) );
  PG_block_79 PG_0_17 ( .A(A[17]), .B(B[17]), .G(\g_vett[0][17] ), .P(
        \p_vett[0][17] ) );
  PG_block_78 PG_0_18 ( .A(A[18]), .B(B[18]), .G(\g_vett[0][18] ), .P(
        \p_vett[0][18] ) );
  PG_block_77 PG_0_19 ( .A(A[19]), .B(B[19]), .G(\g_vett[0][19] ), .P(
        \p_vett[0][19] ) );
  PG_block_76 PG_0_20 ( .A(A[20]), .B(B[20]), .G(\g_vett[0][20] ), .P(
        \p_vett[0][20] ) );
  PG_block_75 PG_0_21 ( .A(A[21]), .B(B[21]), .G(\g_vett[0][21] ), .P(
        \p_vett[0][21] ) );
  PG_block_74 PG_0_22 ( .A(A[22]), .B(B[22]), .G(\g_vett[0][22] ), .P(
        \p_vett[0][22] ) );
  PG_block_73 PG_0_23 ( .A(A[23]), .B(B[23]), .G(\g_vett[0][23] ), .P(
        \p_vett[0][23] ) );
  PG_block_72 PG_0_24 ( .A(A[24]), .B(B[24]), .G(\g_vett[0][24] ), .P(
        \p_vett[0][24] ) );
  PG_block_71 PG_0_25 ( .A(A[25]), .B(B[25]), .G(\g_vett[0][25] ), .P(
        \p_vett[0][25] ) );
  PG_block_70 PG_0_26 ( .A(A[26]), .B(B[26]), .G(\g_vett[0][26] ), .P(
        \p_vett[0][26] ) );
  PG_block_69 PG_0_27 ( .A(A[27]), .B(B[27]), .G(\g_vett[0][27] ), .P(
        \p_vett[0][27] ) );
  PG_block_68 PG_0_28 ( .A(A[28]), .B(B[28]), .G(\g_vett[0][28] ), .P(
        \p_vett[0][28] ) );
  PG_block_67 PG_0_29 ( .A(A[29]), .B(B[29]), .G(\g_vett[0][29] ), .P(
        \p_vett[0][29] ) );
  PG_block_66 PG_0_30 ( .A(A[30]), .B(B[30]), .G(\g_vett[0][30] ), .P(
        \p_vett[0][30] ) );
  PG_block_65 PG_0_31 ( .A(A[31]), .B(B[31]), .G(\g_vett[0][31] ), .P(
        \p_vett[0][31] ) );
  GENERAL_G_29 G_0_0_0 ( .G_in(\g_vett[0][1] ), .P_in(\p_vett[0][1] ), 
        .G_in_prev(\g_vett[0][0] ), .G_out(\g_vett[1][0] ) );
  GENERAL_PG_81 PG_1_0_0 ( .G_in(\g_vett[0][3] ), .P_in(\p_vett[0][3] ), 
        .G_in_prev(\g_vett[0][2] ), .P_in_prev(\p_vett[0][2] ), .G_out(
        \g_vett[1][1] ), .P_out(\p_vett[1][1] ) );
  GENERAL_G_28 G_1_0_0 ( .G_in(\g_vett[1][1] ), .P_in(\p_vett[1][1] ), 
        .G_in_prev(\g_vett[1][0] ), .G_out(Co[1]) );
  GENERAL_PG_80 PG_2_0_1 ( .G_in(\g_vett[0][5] ), .P_in(\p_vett[0][5] ), 
        .G_in_prev(\g_vett[0][4] ), .P_in_prev(\p_vett[0][4] ), .G_out(
        \g_vett[1][2] ), .P_out(\p_vett[1][2] ) );
  GENERAL_PG_79 PG_3_0_1 ( .G_in(\g_vett[0][7] ), .P_in(\p_vett[0][7] ), 
        .G_in_prev(\g_vett[0][6] ), .P_in_prev(\p_vett[0][6] ), .G_out(
        \g_vett[1][3] ), .P_out(\p_vett[1][3] ) );
  GENERAL_PG_78 PG_4_0_1 ( .G_in(\g_vett[1][3] ), .P_in(\p_vett[1][3] ), 
        .G_in_prev(\g_vett[1][2] ), .P_in_prev(\p_vett[1][2] ), .G_out(
        \g_vett[2][1] ), .P_out(\p_vett[2][1] ) );
  GENERAL_PG_77 PG_2_0_2 ( .G_in(\g_vett[0][9] ), .P_in(\p_vett[0][9] ), 
        .G_in_prev(\g_vett[0][8] ), .P_in_prev(\p_vett[0][8] ), .G_out(
        \g_vett[1][4] ), .P_out(\p_vett[1][4] ) );
  GENERAL_PG_76 PG_3_0_2 ( .G_in(\g_vett[0][11] ), .P_in(\p_vett[0][11] ), 
        .G_in_prev(\g_vett[0][10] ), .P_in_prev(\p_vett[0][10] ), .G_out(
        \g_vett[1][5] ), .P_out(\p_vett[1][5] ) );
  GENERAL_PG_75 PG_4_0_2 ( .G_in(\g_vett[1][5] ), .P_in(\p_vett[1][5] ), 
        .G_in_prev(\g_vett[1][4] ), .P_in_prev(\p_vett[1][4] ), .G_out(
        \g_vett[2][2] ), .P_out(\p_vett[2][2] ) );
  GENERAL_PG_74 PG_2_0_3 ( .G_in(\g_vett[0][13] ), .P_in(\p_vett[0][13] ), 
        .G_in_prev(\g_vett[0][12] ), .P_in_prev(\p_vett[0][12] ), .G_out(
        \g_vett[1][6] ), .P_out(\p_vett[1][6] ) );
  GENERAL_PG_73 PG_3_0_3 ( .G_in(\g_vett[0][15] ), .P_in(\p_vett[0][15] ), 
        .G_in_prev(\g_vett[0][14] ), .P_in_prev(\p_vett[0][14] ), .G_out(
        \g_vett[1][7] ), .P_out(\p_vett[1][7] ) );
  GENERAL_PG_72 PG_4_0_3 ( .G_in(\g_vett[1][7] ), .P_in(\p_vett[1][7] ), 
        .G_in_prev(\g_vett[1][6] ), .P_in_prev(\p_vett[1][6] ), .G_out(
        \g_vett[2][3] ), .P_out(\p_vett[2][3] ) );
  GENERAL_PG_71 PG_2_0_4 ( .G_in(\g_vett[0][17] ), .P_in(\p_vett[0][17] ), 
        .G_in_prev(\g_vett[0][16] ), .P_in_prev(\p_vett[0][16] ), .G_out(
        \g_vett[1][8] ), .P_out(\p_vett[1][8] ) );
  GENERAL_PG_70 PG_3_0_4 ( .G_in(\g_vett[0][19] ), .P_in(\p_vett[0][19] ), 
        .G_in_prev(\g_vett[0][18] ), .P_in_prev(\p_vett[0][18] ), .G_out(
        \g_vett[1][9] ), .P_out(\p_vett[1][9] ) );
  GENERAL_PG_69 PG_4_0_4 ( .G_in(\g_vett[1][9] ), .P_in(\p_vett[1][9] ), 
        .G_in_prev(\g_vett[1][8] ), .P_in_prev(\p_vett[1][8] ), .G_out(
        \g_vett[2][4] ), .P_out(\p_vett[2][4] ) );
  GENERAL_PG_68 PG_2_0_5 ( .G_in(\g_vett[0][21] ), .P_in(\p_vett[0][21] ), 
        .G_in_prev(\g_vett[0][20] ), .P_in_prev(\p_vett[0][20] ), .G_out(
        \g_vett[1][10] ), .P_out(\p_vett[1][10] ) );
  GENERAL_PG_67 PG_3_0_5 ( .G_in(\g_vett[0][23] ), .P_in(\p_vett[0][23] ), 
        .G_in_prev(\g_vett[0][22] ), .P_in_prev(\p_vett[0][22] ), .G_out(
        \g_vett[1][11] ), .P_out(\p_vett[1][11] ) );
  GENERAL_PG_66 PG_4_0_5 ( .G_in(\g_vett[1][11] ), .P_in(\p_vett[1][11] ), 
        .G_in_prev(\g_vett[1][10] ), .P_in_prev(\p_vett[1][10] ), .G_out(
        \g_vett[2][5] ), .P_out(\p_vett[2][5] ) );
  GENERAL_PG_65 PG_2_0_6 ( .G_in(\g_vett[0][25] ), .P_in(\p_vett[0][25] ), 
        .G_in_prev(\g_vett[0][24] ), .P_in_prev(\p_vett[0][24] ), .G_out(
        \g_vett[1][12] ), .P_out(\p_vett[1][12] ) );
  GENERAL_PG_64 PG_3_0_6 ( .G_in(\g_vett[0][27] ), .P_in(\p_vett[0][27] ), 
        .G_in_prev(\g_vett[0][26] ), .P_in_prev(\p_vett[0][26] ), .G_out(
        \g_vett[1][13] ), .P_out(\p_vett[1][13] ) );
  GENERAL_PG_63 PG_4_0_6 ( .G_in(\g_vett[1][13] ), .P_in(\p_vett[1][13] ), 
        .G_in_prev(\g_vett[1][12] ), .P_in_prev(\p_vett[1][12] ), .G_out(
        \g_vett[2][6] ), .P_out(\p_vett[2][6] ) );
  GENERAL_PG_62 PG_2_0_7 ( .G_in(\g_vett[0][29] ), .P_in(\p_vett[0][29] ), 
        .G_in_prev(\g_vett[0][28] ), .P_in_prev(\p_vett[0][28] ), .G_out(
        \g_vett[1][14] ), .P_out(\p_vett[1][14] ) );
  GENERAL_PG_61 PG_3_0_7 ( .G_in(\g_vett[0][31] ), .P_in(\p_vett[0][31] ), 
        .G_in_prev(\g_vett[0][30] ), .P_in_prev(\p_vett[0][30] ), .G_out(
        \g_vett[1][15] ), .P_out(\p_vett[1][15] ) );
  GENERAL_PG_60 PG_4_0_7 ( .G_in(\g_vett[1][15] ), .P_in(\p_vett[1][15] ), 
        .G_in_prev(\g_vett[1][14] ), .P_in_prev(\p_vett[1][14] ), .G_out(
        \g_vett[2][7] ), .P_out(\p_vett[2][7] ) );
  GENERAL_G_27 G_2_1_0 ( .G_in(\g_vett[2][1] ), .P_in(\p_vett[2][1] ), 
        .G_in_prev(Co[1]), .G_out(Co[2]) );
  GENERAL_PG_59 PG_5_1_0 ( .G_in(\g_vett[2][3] ), .P_in(\p_vett[2][3] ), 
        .G_in_prev(\g_vett[2][2] ), .P_in_prev(\p_vett[2][2] ), .G_out(
        \g_vett[3][1] ), .P_out(\p_vett[3][1] ) );
  GENERAL_G_26 G_3_1_0 ( .G_in(\g_vett[2][2] ), .P_in(\p_vett[2][2] ), 
        .G_in_prev(Co[2]), .G_out(Co[3]) );
  GENERAL_G_25 G_4_1_0 ( .G_in(\g_vett[3][1] ), .P_in(\p_vett[3][1] ), 
        .G_in_prev(Co[2]), .G_out(Co[4]) );
  GENERAL_PG_58 PG_6_1_1 ( .G_in(\g_vett[2][5] ), .P_in(\p_vett[2][5] ), 
        .G_in_prev(\g_vett[2][4] ), .P_in_prev(\p_vett[2][4] ), .G_out(
        \g_vett[3][2] ), .P_out(\p_vett[3][2] ) );
  GENERAL_PG_57 PG_7_1_1 ( .G_in(\g_vett[2][7] ), .P_in(\p_vett[2][7] ), 
        .G_in_prev(\g_vett[2][6] ), .P_in_prev(\p_vett[2][6] ), .G_out(
        \g_vett[3][3] ), .P_out(\p_vett[3][3] ) );
  GENERAL_PG_56 PG_8_1_1 ( .G_in(\g_vett[2][6] ), .P_in(\p_vett[2][6] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][2] ), .P_out(\p_vett[4][2] ) );
  GENERAL_PG_55 PG_9_1_1 ( .G_in(\g_vett[3][3] ), .P_in(\p_vett[3][3] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][3] ), .P_out(\p_vett[4][3] ) );
  GENERAL_G_24 G_5_2_0 ( .G_in(\g_vett[2][4] ), .P_in(\p_vett[2][4] ), 
        .G_in_prev(Co[4]), .G_out(Co[5]) );
  GENERAL_G_23 G_6_2_1 ( .G_in(\g_vett[3][2] ), .P_in(\p_vett[3][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[6]) );
  GENERAL_G_22 G_7_2_2 ( .G_in(\g_vett[4][2] ), .P_in(\p_vett[4][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[7]) );
  GENERAL_G_21 G_8_2_3 ( .G_in(\g_vett[4][3] ), .P_in(\p_vett[4][3] ), 
        .G_in_prev(Co[4]) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_48 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_192 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_191 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_190 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_189 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_47 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_188 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_187 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_186 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_185 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_48 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U9 ( .A(SEL), .ZN(n13) );
endmodule


module MUX21_GENERIC_NBIT4_47 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U6 ( .A(SEL), .ZN(n13) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_24 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_48 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_47 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_48 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_47 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_46 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_184 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_183 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_182 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_181 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_45 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_180 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_179 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_178 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_177 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_46 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_45 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_23 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_46 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_45 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_46 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_45 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_44 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_176 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_175 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_174 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_173 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_43 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_172 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_171 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_170 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_169 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_44 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_43 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_22 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_44 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_43 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_44 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_43 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_42 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_168 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_167 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_166 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_165 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_41 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_164 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_163 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_162 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_161 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_42 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_41 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_21 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_42 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_41 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_42 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_41 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_40 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_160 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_159 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_158 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_157 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_39 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_156 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_155 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_154 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_153 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_40 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U8 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
endmodule


module MUX21_GENERIC_NBIT4_39 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_20 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_40 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_39 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_40 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_39 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_38 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_152 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_151 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_150 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_149 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_37 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_148 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_147 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_146 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_145 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_38 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_37 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_19 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_38 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_37 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_38 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_37 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_36 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_144 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_143 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_142 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_141 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_35 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_140 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_139 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_138 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_137 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_36 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U6 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U8 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
endmodule


module MUX21_GENERIC_NBIT4_35 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_18 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_36 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_35 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_36 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_35 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_34 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_136 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_135 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_134 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_133 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_33 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_132 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_131 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_130 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_129 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_34 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_33 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_17 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_34 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_33 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_34 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_33 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module SUMGEN_NBIT32_NBLOCKS8_3 ( A, B, cin_vect, Co, SUM );
  input [31:0] A;
  input [31:0] B;
  input [7:0] cin_vect;
  output [31:0] SUM;
  output Co;


  CSblock_NBIT4_24 block_i_0 ( .A(A[3:0]), .B(B[3:0]), .cin(cin_vect[0]), .Y(
        SUM[3:0]) );
  CSblock_NBIT4_23 block_i_1 ( .A(A[7:4]), .B(B[7:4]), .cin(cin_vect[1]), .Y(
        SUM[7:4]) );
  CSblock_NBIT4_22 block_i_2 ( .A(A[11:8]), .B(B[11:8]), .cin(cin_vect[2]), 
        .Y(SUM[11:8]) );
  CSblock_NBIT4_21 block_i_3 ( .A(A[15:12]), .B(B[15:12]), .cin(cin_vect[3]), 
        .Y(SUM[15:12]) );
  CSblock_NBIT4_20 block_i_4 ( .A(A[19:16]), .B(B[19:16]), .cin(cin_vect[4]), 
        .Y(SUM[19:16]) );
  CSblock_NBIT4_19 block_i_5 ( .A(A[23:20]), .B(B[23:20]), .cin(cin_vect[5]), 
        .Y(SUM[23:20]) );
  CSblock_NBIT4_18 block_i_6 ( .A(A[27:24]), .B(B[27:24]), .cin(cin_vect[6]), 
        .Y(SUM[27:24]) );
  CSblock_NBIT4_17 block_i_7 ( .A(A[31:28]), .B(B[31:28]), .cin(cin_vect[7]), 
        .Y(SUM[31:28]), .Co(Co) );
endmodule


module P4_ADDER_NBIT32_NBIT_PER_BLOCK4_3 ( A, B, Cin, Cout, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input Cin;
  output Cout;

  wire   [7:0] outCarryGen;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 CG ( .A(A), .B(B), .Cin(Cin), .Co(
        outCarryGen) );
  SUMGEN_NBIT32_NBLOCKS8_3 SG ( .A(A), .B(B), .cin_vect(outCarryGen), .Co(Cout), .SUM(Y) );
endmodule


module PG_block_64 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_20 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module PG_block_63 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_62 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_61 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_60 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_59 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_58 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_57 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_56 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_55 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_54 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_53 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_52 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_51 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_50 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_49 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_48 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_47 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_46 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_45 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_44 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_43 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_42 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_41 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_40 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_39 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_38 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_37 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_36 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_35 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_34 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_block_33 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GENERAL_G_19 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_54 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_18 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_53 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_52 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_51 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_50 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_49 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_48 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_47 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_46 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_45 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_44 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_43 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_42 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_41 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_40 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_39 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_38 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_37 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_36 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_35 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_34 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_33 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_G_17 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_32 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_16 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_15 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_31 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
  AND2_X1 U3 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
endmodule


module GENERAL_PG_30 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_29 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  AND2_X1 U1 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  INV_X1 U2 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_PG_28 ( G_in, P_in, G_in_prev, P_in_prev, G_out, P_out );
  input G_in, P_in, G_in_prev, P_in_prev;
  output G_out, P_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AND2_X1 U2 ( .A1(P_in_prev), .A2(P_in), .ZN(P_out) );
  AOI21_X1 U3 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_14 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_13 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_12 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module GENERAL_G_11 ( G_in, P_in, G_in_prev, G_out );
  input G_in, P_in, G_in_prev;
  output G_out;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(G_out) );
  AOI21_X1 U2 ( .B1(P_in), .B2(G_in_prev), .A(G_in), .ZN(n4) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   Cin, first_generate, \p_vett[4][3] , \p_vett[4][2] , \p_vett[3][3] ,
         \p_vett[3][2] , \p_vett[3][1] , \p_vett[2][7] , \p_vett[2][6] ,
         \p_vett[2][5] , \p_vett[2][4] , \p_vett[2][3] , \p_vett[2][2] ,
         \p_vett[2][1] , \p_vett[1][15] , \p_vett[1][14] , \p_vett[1][13] ,
         \p_vett[1][12] , \p_vett[1][11] , \p_vett[1][10] , \p_vett[1][9] ,
         \p_vett[1][8] , \p_vett[1][7] , \p_vett[1][6] , \p_vett[1][5] ,
         \p_vett[1][4] , \p_vett[1][3] , \p_vett[1][2] , \p_vett[1][1] ,
         \p_vett[0][31] , \p_vett[0][30] , \p_vett[0][29] , \p_vett[0][28] ,
         \p_vett[0][27] , \p_vett[0][26] , \p_vett[0][25] , \p_vett[0][24] ,
         \p_vett[0][23] , \p_vett[0][22] , \p_vett[0][21] , \p_vett[0][20] ,
         \p_vett[0][19] , \p_vett[0][18] , \p_vett[0][17] , \p_vett[0][16] ,
         \p_vett[0][15] , \p_vett[0][14] , \p_vett[0][13] , \p_vett[0][12] ,
         \p_vett[0][11] , \p_vett[0][10] , \p_vett[0][9] , \p_vett[0][8] ,
         \p_vett[0][7] , \p_vett[0][6] , \p_vett[0][5] , \p_vett[0][4] ,
         \p_vett[0][3] , \p_vett[0][2] , \p_vett[0][1] , \p_vett[0][0] ,
         \g_vett[4][3] , \g_vett[4][2] , \g_vett[3][3] , \g_vett[3][2] ,
         \g_vett[3][1] , \g_vett[2][7] , \g_vett[2][6] , \g_vett[2][5] ,
         \g_vett[2][4] , \g_vett[2][3] , \g_vett[2][2] , \g_vett[2][1] ,
         \g_vett[1][15] , \g_vett[1][14] , \g_vett[1][13] , \g_vett[1][12] ,
         \g_vett[1][11] , \g_vett[1][10] , \g_vett[1][9] , \g_vett[1][8] ,
         \g_vett[1][7] , \g_vett[1][6] , \g_vett[1][5] , \g_vett[1][4] ,
         \g_vett[1][3] , \g_vett[1][2] , \g_vett[1][1] , \g_vett[1][0] ,
         \g_vett[0][31] , \g_vett[0][30] , \g_vett[0][29] , \g_vett[0][28] ,
         \g_vett[0][27] , \g_vett[0][26] , \g_vett[0][25] , \g_vett[0][24] ,
         \g_vett[0][23] , \g_vett[0][22] , \g_vett[0][21] , \g_vett[0][20] ,
         \g_vett[0][19] , \g_vett[0][18] , \g_vett[0][17] , \g_vett[0][16] ,
         \g_vett[0][15] , \g_vett[0][14] , \g_vett[0][13] , \g_vett[0][12] ,
         \g_vett[0][11] , \g_vett[0][10] , \g_vett[0][9] , \g_vett[0][8] ,
         \g_vett[0][7] , \g_vett[0][6] , \g_vett[0][5] , \g_vett[0][4] ,
         \g_vett[0][3] , \g_vett[0][2] , \g_vett[0][1] , \g_vett[0][0] ;
  assign Co[0] = Cin;

  PG_block_64 PGblock_first ( .A(A[0]), .B(B[0]), .G(first_generate), .P(
        \p_vett[0][0] ) );
  GENERAL_G_20 G_first ( .G_in(first_generate), .P_in(\p_vett[0][0] ), 
        .G_in_prev(Cin), .G_out(\g_vett[0][0] ) );
  PG_block_63 PG_0_1 ( .A(A[1]), .B(B[1]), .G(\g_vett[0][1] ), .P(
        \p_vett[0][1] ) );
  PG_block_62 PG_0_2 ( .A(A[2]), .B(B[2]), .G(\g_vett[0][2] ), .P(
        \p_vett[0][2] ) );
  PG_block_61 PG_0_3 ( .A(A[3]), .B(B[3]), .G(\g_vett[0][3] ), .P(
        \p_vett[0][3] ) );
  PG_block_60 PG_0_4 ( .A(A[4]), .B(B[4]), .G(\g_vett[0][4] ), .P(
        \p_vett[0][4] ) );
  PG_block_59 PG_0_5 ( .A(A[5]), .B(B[5]), .G(\g_vett[0][5] ), .P(
        \p_vett[0][5] ) );
  PG_block_58 PG_0_6 ( .A(A[6]), .B(B[6]), .G(\g_vett[0][6] ), .P(
        \p_vett[0][6] ) );
  PG_block_57 PG_0_7 ( .A(A[7]), .B(B[7]), .G(\g_vett[0][7] ), .P(
        \p_vett[0][7] ) );
  PG_block_56 PG_0_8 ( .A(A[8]), .B(B[8]), .G(\g_vett[0][8] ), .P(
        \p_vett[0][8] ) );
  PG_block_55 PG_0_9 ( .A(A[9]), .B(B[9]), .G(\g_vett[0][9] ), .P(
        \p_vett[0][9] ) );
  PG_block_54 PG_0_10 ( .A(A[10]), .B(B[10]), .G(\g_vett[0][10] ), .P(
        \p_vett[0][10] ) );
  PG_block_53 PG_0_11 ( .A(A[11]), .B(B[11]), .G(\g_vett[0][11] ), .P(
        \p_vett[0][11] ) );
  PG_block_52 PG_0_12 ( .A(A[12]), .B(B[12]), .G(\g_vett[0][12] ), .P(
        \p_vett[0][12] ) );
  PG_block_51 PG_0_13 ( .A(A[13]), .B(B[13]), .G(\g_vett[0][13] ), .P(
        \p_vett[0][13] ) );
  PG_block_50 PG_0_14 ( .A(A[14]), .B(B[14]), .G(\g_vett[0][14] ), .P(
        \p_vett[0][14] ) );
  PG_block_49 PG_0_15 ( .A(A[15]), .B(B[15]), .G(\g_vett[0][15] ), .P(
        \p_vett[0][15] ) );
  PG_block_48 PG_0_16 ( .A(A[16]), .B(B[16]), .G(\g_vett[0][16] ), .P(
        \p_vett[0][16] ) );
  PG_block_47 PG_0_17 ( .A(A[17]), .B(B[17]), .G(\g_vett[0][17] ), .P(
        \p_vett[0][17] ) );
  PG_block_46 PG_0_18 ( .A(A[18]), .B(B[18]), .G(\g_vett[0][18] ), .P(
        \p_vett[0][18] ) );
  PG_block_45 PG_0_19 ( .A(A[19]), .B(B[19]), .G(\g_vett[0][19] ), .P(
        \p_vett[0][19] ) );
  PG_block_44 PG_0_20 ( .A(A[20]), .B(B[20]), .G(\g_vett[0][20] ), .P(
        \p_vett[0][20] ) );
  PG_block_43 PG_0_21 ( .A(A[21]), .B(B[21]), .G(\g_vett[0][21] ), .P(
        \p_vett[0][21] ) );
  PG_block_42 PG_0_22 ( .A(A[22]), .B(B[22]), .G(\g_vett[0][22] ), .P(
        \p_vett[0][22] ) );
  PG_block_41 PG_0_23 ( .A(A[23]), .B(B[23]), .G(\g_vett[0][23] ), .P(
        \p_vett[0][23] ) );
  PG_block_40 PG_0_24 ( .A(A[24]), .B(B[24]), .G(\g_vett[0][24] ), .P(
        \p_vett[0][24] ) );
  PG_block_39 PG_0_25 ( .A(A[25]), .B(B[25]), .G(\g_vett[0][25] ), .P(
        \p_vett[0][25] ) );
  PG_block_38 PG_0_26 ( .A(A[26]), .B(B[26]), .G(\g_vett[0][26] ), .P(
        \p_vett[0][26] ) );
  PG_block_37 PG_0_27 ( .A(A[27]), .B(B[27]), .G(\g_vett[0][27] ), .P(
        \p_vett[0][27] ) );
  PG_block_36 PG_0_28 ( .A(A[28]), .B(B[28]), .G(\g_vett[0][28] ), .P(
        \p_vett[0][28] ) );
  PG_block_35 PG_0_29 ( .A(A[29]), .B(B[29]), .G(\g_vett[0][29] ), .P(
        \p_vett[0][29] ) );
  PG_block_34 PG_0_30 ( .A(A[30]), .B(B[30]), .G(\g_vett[0][30] ), .P(
        \p_vett[0][30] ) );
  PG_block_33 PG_0_31 ( .A(A[31]), .B(B[31]), .G(\g_vett[0][31] ), .P(
        \p_vett[0][31] ) );
  GENERAL_G_19 G_0_0_0 ( .G_in(\g_vett[0][1] ), .P_in(\p_vett[0][1] ), 
        .G_in_prev(\g_vett[0][0] ), .G_out(\g_vett[1][0] ) );
  GENERAL_PG_54 PG_1_0_0 ( .G_in(\g_vett[0][3] ), .P_in(\p_vett[0][3] ), 
        .G_in_prev(\g_vett[0][2] ), .P_in_prev(\p_vett[0][2] ), .G_out(
        \g_vett[1][1] ), .P_out(\p_vett[1][1] ) );
  GENERAL_G_18 G_1_0_0 ( .G_in(\g_vett[1][1] ), .P_in(\p_vett[1][1] ), 
        .G_in_prev(\g_vett[1][0] ), .G_out(Co[1]) );
  GENERAL_PG_53 PG_2_0_1 ( .G_in(\g_vett[0][5] ), .P_in(\p_vett[0][5] ), 
        .G_in_prev(\g_vett[0][4] ), .P_in_prev(\p_vett[0][4] ), .G_out(
        \g_vett[1][2] ), .P_out(\p_vett[1][2] ) );
  GENERAL_PG_52 PG_3_0_1 ( .G_in(\g_vett[0][7] ), .P_in(\p_vett[0][7] ), 
        .G_in_prev(\g_vett[0][6] ), .P_in_prev(\p_vett[0][6] ), .G_out(
        \g_vett[1][3] ), .P_out(\p_vett[1][3] ) );
  GENERAL_PG_51 PG_4_0_1 ( .G_in(\g_vett[1][3] ), .P_in(\p_vett[1][3] ), 
        .G_in_prev(\g_vett[1][2] ), .P_in_prev(\p_vett[1][2] ), .G_out(
        \g_vett[2][1] ), .P_out(\p_vett[2][1] ) );
  GENERAL_PG_50 PG_2_0_2 ( .G_in(\g_vett[0][9] ), .P_in(\p_vett[0][9] ), 
        .G_in_prev(\g_vett[0][8] ), .P_in_prev(\p_vett[0][8] ), .G_out(
        \g_vett[1][4] ), .P_out(\p_vett[1][4] ) );
  GENERAL_PG_49 PG_3_0_2 ( .G_in(\g_vett[0][11] ), .P_in(\p_vett[0][11] ), 
        .G_in_prev(\g_vett[0][10] ), .P_in_prev(\p_vett[0][10] ), .G_out(
        \g_vett[1][5] ), .P_out(\p_vett[1][5] ) );
  GENERAL_PG_48 PG_4_0_2 ( .G_in(\g_vett[1][5] ), .P_in(\p_vett[1][5] ), 
        .G_in_prev(\g_vett[1][4] ), .P_in_prev(\p_vett[1][4] ), .G_out(
        \g_vett[2][2] ), .P_out(\p_vett[2][2] ) );
  GENERAL_PG_47 PG_2_0_3 ( .G_in(\g_vett[0][13] ), .P_in(\p_vett[0][13] ), 
        .G_in_prev(\g_vett[0][12] ), .P_in_prev(\p_vett[0][12] ), .G_out(
        \g_vett[1][6] ), .P_out(\p_vett[1][6] ) );
  GENERAL_PG_46 PG_3_0_3 ( .G_in(\g_vett[0][15] ), .P_in(\p_vett[0][15] ), 
        .G_in_prev(\g_vett[0][14] ), .P_in_prev(\p_vett[0][14] ), .G_out(
        \g_vett[1][7] ), .P_out(\p_vett[1][7] ) );
  GENERAL_PG_45 PG_4_0_3 ( .G_in(\g_vett[1][7] ), .P_in(\p_vett[1][7] ), 
        .G_in_prev(\g_vett[1][6] ), .P_in_prev(\p_vett[1][6] ), .G_out(
        \g_vett[2][3] ), .P_out(\p_vett[2][3] ) );
  GENERAL_PG_44 PG_2_0_4 ( .G_in(\g_vett[0][17] ), .P_in(\p_vett[0][17] ), 
        .G_in_prev(\g_vett[0][16] ), .P_in_prev(\p_vett[0][16] ), .G_out(
        \g_vett[1][8] ), .P_out(\p_vett[1][8] ) );
  GENERAL_PG_43 PG_3_0_4 ( .G_in(\g_vett[0][19] ), .P_in(\p_vett[0][19] ), 
        .G_in_prev(\g_vett[0][18] ), .P_in_prev(\p_vett[0][18] ), .G_out(
        \g_vett[1][9] ), .P_out(\p_vett[1][9] ) );
  GENERAL_PG_42 PG_4_0_4 ( .G_in(\g_vett[1][9] ), .P_in(\p_vett[1][9] ), 
        .G_in_prev(\g_vett[1][8] ), .P_in_prev(\p_vett[1][8] ), .G_out(
        \g_vett[2][4] ), .P_out(\p_vett[2][4] ) );
  GENERAL_PG_41 PG_2_0_5 ( .G_in(\g_vett[0][21] ), .P_in(\p_vett[0][21] ), 
        .G_in_prev(\g_vett[0][20] ), .P_in_prev(\p_vett[0][20] ), .G_out(
        \g_vett[1][10] ), .P_out(\p_vett[1][10] ) );
  GENERAL_PG_40 PG_3_0_5 ( .G_in(\g_vett[0][23] ), .P_in(\p_vett[0][23] ), 
        .G_in_prev(\g_vett[0][22] ), .P_in_prev(\p_vett[0][22] ), .G_out(
        \g_vett[1][11] ), .P_out(\p_vett[1][11] ) );
  GENERAL_PG_39 PG_4_0_5 ( .G_in(\g_vett[1][11] ), .P_in(\p_vett[1][11] ), 
        .G_in_prev(\g_vett[1][10] ), .P_in_prev(\p_vett[1][10] ), .G_out(
        \g_vett[2][5] ), .P_out(\p_vett[2][5] ) );
  GENERAL_PG_38 PG_2_0_6 ( .G_in(\g_vett[0][25] ), .P_in(\p_vett[0][25] ), 
        .G_in_prev(\g_vett[0][24] ), .P_in_prev(\p_vett[0][24] ), .G_out(
        \g_vett[1][12] ), .P_out(\p_vett[1][12] ) );
  GENERAL_PG_37 PG_3_0_6 ( .G_in(\g_vett[0][27] ), .P_in(\p_vett[0][27] ), 
        .G_in_prev(\g_vett[0][26] ), .P_in_prev(\p_vett[0][26] ), .G_out(
        \g_vett[1][13] ), .P_out(\p_vett[1][13] ) );
  GENERAL_PG_36 PG_4_0_6 ( .G_in(\g_vett[1][13] ), .P_in(\p_vett[1][13] ), 
        .G_in_prev(\g_vett[1][12] ), .P_in_prev(\p_vett[1][12] ), .G_out(
        \g_vett[2][6] ), .P_out(\p_vett[2][6] ) );
  GENERAL_PG_35 PG_2_0_7 ( .G_in(\g_vett[0][29] ), .P_in(\p_vett[0][29] ), 
        .G_in_prev(\g_vett[0][28] ), .P_in_prev(\p_vett[0][28] ), .G_out(
        \g_vett[1][14] ), .P_out(\p_vett[1][14] ) );
  GENERAL_PG_34 PG_3_0_7 ( .G_in(\g_vett[0][31] ), .P_in(\p_vett[0][31] ), 
        .G_in_prev(\g_vett[0][30] ), .P_in_prev(\p_vett[0][30] ), .G_out(
        \g_vett[1][15] ), .P_out(\p_vett[1][15] ) );
  GENERAL_PG_33 PG_4_0_7 ( .G_in(\g_vett[1][15] ), .P_in(\p_vett[1][15] ), 
        .G_in_prev(\g_vett[1][14] ), .P_in_prev(\p_vett[1][14] ), .G_out(
        \g_vett[2][7] ), .P_out(\p_vett[2][7] ) );
  GENERAL_G_17 G_2_1_0 ( .G_in(\g_vett[2][1] ), .P_in(\p_vett[2][1] ), 
        .G_in_prev(Co[1]), .G_out(Co[2]) );
  GENERAL_PG_32 PG_5_1_0 ( .G_in(\g_vett[2][3] ), .P_in(\p_vett[2][3] ), 
        .G_in_prev(\g_vett[2][2] ), .P_in_prev(\p_vett[2][2] ), .G_out(
        \g_vett[3][1] ), .P_out(\p_vett[3][1] ) );
  GENERAL_G_16 G_3_1_0 ( .G_in(\g_vett[2][2] ), .P_in(\p_vett[2][2] ), 
        .G_in_prev(Co[2]), .G_out(Co[3]) );
  GENERAL_G_15 G_4_1_0 ( .G_in(\g_vett[3][1] ), .P_in(\p_vett[3][1] ), 
        .G_in_prev(Co[2]), .G_out(Co[4]) );
  GENERAL_PG_31 PG_6_1_1 ( .G_in(\g_vett[2][5] ), .P_in(\p_vett[2][5] ), 
        .G_in_prev(\g_vett[2][4] ), .P_in_prev(\p_vett[2][4] ), .G_out(
        \g_vett[3][2] ), .P_out(\p_vett[3][2] ) );
  GENERAL_PG_30 PG_7_1_1 ( .G_in(\g_vett[2][7] ), .P_in(\p_vett[2][7] ), 
        .G_in_prev(\g_vett[2][6] ), .P_in_prev(\p_vett[2][6] ), .G_out(
        \g_vett[3][3] ), .P_out(\p_vett[3][3] ) );
  GENERAL_PG_29 PG_8_1_1 ( .G_in(\g_vett[2][6] ), .P_in(\p_vett[2][6] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][2] ), .P_out(\p_vett[4][2] ) );
  GENERAL_PG_28 PG_9_1_1 ( .G_in(\g_vett[3][3] ), .P_in(\p_vett[3][3] ), 
        .G_in_prev(\g_vett[3][2] ), .P_in_prev(\p_vett[3][2] ), .G_out(
        \g_vett[4][3] ), .P_out(\p_vett[4][3] ) );
  GENERAL_G_14 G_5_2_0 ( .G_in(\g_vett[2][4] ), .P_in(\p_vett[2][4] ), 
        .G_in_prev(Co[4]), .G_out(Co[5]) );
  GENERAL_G_13 G_6_2_1 ( .G_in(\g_vett[3][2] ), .P_in(\p_vett[3][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[6]) );
  GENERAL_G_12 G_7_2_2 ( .G_in(\g_vett[4][2] ), .P_in(\p_vett[4][2] ), 
        .G_in_prev(Co[4]), .G_out(Co[7]) );
  GENERAL_G_11 G_8_2_3 ( .G_in(\g_vett[4][3] ), .P_in(\p_vett[4][3] ), 
        .G_in_prev(Co[4]) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_32 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_128 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_127 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_126 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_125 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_31 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_124 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_123 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_122 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_121 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_32 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U2 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U9 ( .A(SEL), .ZN(n13) );
endmodule


module MUX21_GENERIC_NBIT4_31 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U6 ( .A(SEL), .ZN(n13) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_16 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_32 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_31 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_32 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_31 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_120 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_119 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_118 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_117 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_116 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_115 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_114 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_113 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_30 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_29 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_15 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_30 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_29 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_30 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_29 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_112 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_111 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_110 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_109 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_108 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_107 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_106 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_105 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_28 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_27 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_14 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_28 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_27 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_28 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_27 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_104 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_103 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_102 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_101 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_100 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_99 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_98 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_97 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_26 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_25 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_13 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_26 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_25 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_26 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_25 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_96 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_95 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_94 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_93 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_92 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_91 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_90 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_89 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_24 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
  INV_X1 U4 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U6 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U8 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
endmodule


module MUX21_GENERIC_NBIT4_23 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_12 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_24 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_23 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_24 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_23 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_88 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_87 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_86 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_85 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_84 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_83 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_82 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_81 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_22 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_21 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_11 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_22 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_21 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_22 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_21 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_80 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_79 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_78 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_77 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_76 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_75 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_74 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_73 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_20 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_19 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_10 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_20 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_19 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_20 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_19 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module RCA_NBIT4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_72 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_71 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_70 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_69 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_NBIT4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_68 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_67 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_66 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_65 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_NBIT4_18 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  AOI22_X1 U3 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  INV_X1 U4 ( .A(n15), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(Y[2]) );
  AOI22_X1 U7 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module MUX21_GENERIC_NBIT4_17 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n15), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n16), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n17), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(A[0]), .A2(n13), .B1(B[0]), .B2(SEL), .ZN(n14) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n13), .B1(B[1]), .B2(SEL), .ZN(n15) );
  AOI22_X1 U8 ( .A1(A[2]), .A2(n13), .B1(B[2]), .B2(SEL), .ZN(n16) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n13), .B1(SEL), .B2(B[3]), .ZN(n17) );
endmodule


module CSblock_NBIT4_9 ( A, B, cin, Y, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input cin;
  output Co;
  wire   \cout0[0] , \cout1[0] ;
  wire   [3:0] out0;
  wire   [3:0] out1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  RCA_NBIT4_18 add0 ( .A(A), .B(B), .Ci(1'b0), .S(out0), .Co(\cout0[0] ) );
  RCA_NBIT4_17 add1 ( .A(A), .B(B), .Ci(1'b0), .S(out1), .Co(\cout1[0] ) );
  MUX21_GENERIC_NBIT4_18 muxSum ( .A(out0), .B(out1), .SEL(cin), .Y(Y) );
  MUX21_GENERIC_NBIT4_17 muxCout ( .A({1'b0, 1'b0, 1'b0, \cout0[0] }), .B({
        1'b0, 1'b0, 1'b0, \cout1[0] }), .SEL(cin), .Y({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, Co}) );
endmodule


module SUMGEN_NBIT32_NBLOCKS8_2 ( A, B, cin_vect, Co, SUM );
  input [31:0] A;
  input [31:0] B;
  input [7:0] cin_vect;
  output [31:0] SUM;
  output Co;


  CSblock_NBIT4_16 block_i_0 ( .A(A[3:0]), .B(B[3:0]), .cin(cin_vect[0]), .Y(
        SUM[3:0]) );
  CSblock_NBIT4_15 block_i_1 ( .A(A[7:4]), .B(B[7:4]), .cin(cin_vect[1]), .Y(
        SUM[7:4]) );
  CSblock_NBIT4_14 block_i_2 ( .A(A[11:8]), .B(B[11:8]), .cin(cin_vect[2]), 
        .Y(SUM[11:8]) );
  CSblock_NBIT4_13 block_i_3 ( .A(A[15:12]), .B(B[15:12]), .cin(cin_vect[3]), 
        .Y(SUM[15:12]) );
  CSblock_NBIT4_12 block_i_4 ( .A(A[19:16]), .B(B[19:16]), .cin(cin_vect[4]), 
        .Y(SUM[19:16]) );
  CSblock_NBIT4_11 block_i_5 ( .A(A[23:20]), .B(B[23:20]), .cin(cin_vect[5]), 
        .Y(SUM[23:20]) );
  CSblock_NBIT4_10 block_i_6 ( .A(A[27:24]), .B(B[27:24]), .cin(cin_vect[6]), 
        .Y(SUM[27:24]) );
  CSblock_NBIT4_9 block_i_7 ( .A(A[31:28]), .B(B[31:28]), .cin(cin_vect[7]), 
        .Y(SUM[31:28]), .Co(Co) );
endmodule


module P4_ADDER_NBIT32_NBIT_PER_BLOCK4_2 ( A, B, Cin, Cout, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input Cin;
  output Cout;

  wire   [7:0] outCarryGen;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 CG ( .A(A), .B(B), .Cin(Cin), .Co(
        outCarryGen) );
  SUMGEN_NBIT32_NBLOCKS8_2 SG ( .A(A), .B(B), .cin_vect(outCarryGen), .Co(Cout), .SUM(Y) );
endmodule


module REG_GEN_NBIT32_7 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n50), .Q(Q[31]), .QN(n148) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n50), .Q(Q[30]), .QN(n147) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n50), .Q(Q[29]), .QN(n146) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n50), .Q(Q[28]), .QN(n145) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n50), .Q(Q[27]), .QN(n144) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n50), .Q(Q[26]), .QN(n143) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n50), .Q(Q[25]), .QN(n142) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n50), .Q(Q[24]), .QN(n141) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n50), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n50), .Q(Q[22]), .QN(n139) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n50), .Q(Q[21]), .QN(n138) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n50), .Q(Q[20]), .QN(n137) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n136) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n135) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n51), .Q(Q[17]), .QN(n134) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n133) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n132) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n131) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n51), .Q(Q[13]), .QN(n130) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n51), .Q(Q[12]), .QN(n129) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n51), .Q(Q[11]), .QN(n128) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n51), .Q(Q[10]), .QN(n127) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n51), .Q(Q[9]), .QN(n126) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n51), .Q(Q[8]), .QN(n125) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n52), .Q(Q[7]), .QN(n124) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n52), .Q(Q[6]), .QN(n123) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n52), .Q(Q[5]), .QN(n122) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n52), .Q(Q[4]), .QN(n121) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n52), .Q(Q[3]), .QN(n120) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n52), .Q(Q[2]), .QN(n119) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n52), .Q(Q[1]), .QN(n118) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n52), .Q(Q[0]), .QN(n117) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n44) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n136), .A2(n39), .B1(n47), .B2(n101), .ZN(n16) );
  INV_X1 U20 ( .A(D[19]), .ZN(n101) );
  OAI22_X1 U21 ( .A1(n129), .A2(n40), .B1(n45), .B2(n100), .ZN(n23) );
  INV_X1 U22 ( .A(D[12]), .ZN(n100) );
  OAI22_X1 U23 ( .A1(n130), .A2(n40), .B1(n45), .B2(n99), .ZN(n22) );
  INV_X1 U24 ( .A(D[13]), .ZN(n99) );
  OAI22_X1 U25 ( .A1(n131), .A2(n39), .B1(n46), .B2(n98), .ZN(n21) );
  INV_X1 U26 ( .A(D[14]), .ZN(n98) );
  OAI22_X1 U27 ( .A1(n143), .A2(n40), .B1(n41), .B2(n110), .ZN(n9) );
  INV_X1 U28 ( .A(D[26]), .ZN(n110) );
  OAI22_X1 U29 ( .A1(n144), .A2(n39), .B1(n41), .B2(n109), .ZN(n8) );
  INV_X1 U30 ( .A(D[27]), .ZN(n109) );
  OAI22_X1 U31 ( .A1(n145), .A2(n40), .B1(n41), .B2(n116), .ZN(n7) );
  INV_X1 U32 ( .A(D[28]), .ZN(n116) );
  OAI22_X1 U33 ( .A1(n146), .A2(n39), .B1(n41), .B2(n115), .ZN(n6) );
  INV_X1 U34 ( .A(D[29]), .ZN(n115) );
  OAI22_X1 U35 ( .A1(n147), .A2(n40), .B1(n42), .B2(n114), .ZN(n5) );
  INV_X1 U36 ( .A(D[30]), .ZN(n114) );
  OAI22_X1 U37 ( .A1(n148), .A2(n39), .B1(n42), .B2(n113), .ZN(n4) );
  INV_X1 U38 ( .A(D[31]), .ZN(n113) );
  OAI22_X1 U39 ( .A1(n132), .A2(n39), .B1(n46), .B2(n65), .ZN(n20) );
  INV_X1 U40 ( .A(D[15]), .ZN(n65) );
  OAI22_X1 U41 ( .A1(n133), .A2(n39), .B1(n46), .B2(n104), .ZN(n19) );
  INV_X1 U42 ( .A(D[16]), .ZN(n104) );
  OAI22_X1 U43 ( .A1(n134), .A2(n39), .B1(n46), .B2(n103), .ZN(n18) );
  INV_X1 U44 ( .A(D[17]), .ZN(n103) );
  OAI22_X1 U45 ( .A1(n135), .A2(n39), .B1(n47), .B2(n102), .ZN(n17) );
  INV_X1 U46 ( .A(D[18]), .ZN(n102) );
  OAI22_X1 U47 ( .A1(n137), .A2(n39), .B1(n47), .B2(n108), .ZN(n15) );
  INV_X1 U48 ( .A(D[20]), .ZN(n108) );
  OAI22_X1 U49 ( .A1(n138), .A2(n39), .B1(n47), .B2(n107), .ZN(n14) );
  INV_X1 U50 ( .A(D[21]), .ZN(n107) );
  OAI22_X1 U51 ( .A1(n139), .A2(n39), .B1(n48), .B2(n106), .ZN(n13) );
  INV_X1 U52 ( .A(D[22]), .ZN(n106) );
  OAI22_X1 U53 ( .A1(n140), .A2(n39), .B1(n48), .B2(n105), .ZN(n12) );
  INV_X1 U54 ( .A(D[23]), .ZN(n105) );
  OAI22_X1 U55 ( .A1(n141), .A2(n39), .B1(n48), .B2(n112), .ZN(n11) );
  INV_X1 U56 ( .A(D[24]), .ZN(n112) );
  OAI22_X1 U57 ( .A1(n142), .A2(n39), .B1(n48), .B2(n111), .ZN(n10) );
  INV_X1 U58 ( .A(D[25]), .ZN(n111) );
  OAI22_X1 U59 ( .A1(n117), .A2(n40), .B1(n42), .B2(n56), .ZN(n35) );
  INV_X1 U60 ( .A(D[0]), .ZN(n56) );
  OAI22_X1 U61 ( .A1(n125), .A2(n40), .B1(n44), .B2(n64), .ZN(n27) );
  INV_X1 U62 ( .A(D[8]), .ZN(n64) );
  OAI22_X1 U63 ( .A1(n126), .A2(n40), .B1(n44), .B2(n63), .ZN(n26) );
  INV_X1 U64 ( .A(D[9]), .ZN(n63) );
  OAI22_X1 U65 ( .A1(n127), .A2(n40), .B1(n45), .B2(n62), .ZN(n25) );
  INV_X1 U66 ( .A(D[10]), .ZN(n62) );
  OAI22_X1 U67 ( .A1(n121), .A2(n40), .B1(n43), .B2(n60), .ZN(n31) );
  INV_X1 U68 ( .A(D[4]), .ZN(n60) );
  OAI22_X1 U69 ( .A1(n122), .A2(n40), .B1(n43), .B2(n59), .ZN(n30) );
  INV_X1 U70 ( .A(D[5]), .ZN(n59) );
  OAI22_X1 U71 ( .A1(n123), .A2(n40), .B1(n44), .B2(n58), .ZN(n29) );
  INV_X1 U72 ( .A(D[6]), .ZN(n58) );
  OAI22_X1 U73 ( .A1(n128), .A2(n40), .B1(n45), .B2(n61), .ZN(n24) );
  INV_X1 U74 ( .A(D[11]), .ZN(n61) );
  OAI22_X1 U75 ( .A1(n124), .A2(n40), .B1(n44), .B2(n57), .ZN(n28) );
  INV_X1 U76 ( .A(D[7]), .ZN(n57) );
  OAI22_X1 U77 ( .A1(n118), .A2(n39), .B1(n42), .B2(n55), .ZN(n34) );
  INV_X1 U78 ( .A(D[1]), .ZN(n55) );
  OAI22_X1 U79 ( .A1(n119), .A2(n40), .B1(n43), .B2(n54), .ZN(n33) );
  INV_X1 U80 ( .A(D[2]), .ZN(n54) );
  OAI22_X1 U81 ( .A1(n120), .A2(n40), .B1(n43), .B2(n53), .ZN(n32) );
  INV_X1 U82 ( .A(D[3]), .ZN(n53) );
endmodule


module REG_GEN_NBIT32_6 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n50), .Q(Q[31]), .QN(n148) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n50), .Q(Q[30]), .QN(n147) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n50), .Q(Q[29]), .QN(n146) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n50), .Q(Q[28]), .QN(n145) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n50), .Q(Q[27]), .QN(n144) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n50), .Q(Q[26]), .QN(n143) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n50), .Q(Q[25]), .QN(n142) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n50), .Q(Q[24]), .QN(n141) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n50), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n50), .Q(Q[22]), .QN(n139) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n50), .Q(Q[21]), .QN(n138) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n50), .Q(Q[20]), .QN(n137) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n136) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n135) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n51), .Q(Q[17]), .QN(n134) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n133) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n132) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n131) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n51), .Q(Q[13]), .QN(n130) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n51), .Q(Q[12]), .QN(n129) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n51), .Q(Q[11]), .QN(n128) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n51), .Q(Q[10]), .QN(n127) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n51), .Q(Q[9]), .QN(n126) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n51), .Q(Q[8]), .QN(n125) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n52), .Q(Q[7]), .QN(n124) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n52), .Q(Q[6]), .QN(n123) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n52), .Q(Q[5]), .QN(n122) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n52), .Q(Q[4]), .QN(n121) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n52), .Q(Q[3]), .QN(n120) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n52), .Q(Q[2]), .QN(n119) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n52), .Q(Q[1]), .QN(n118) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n52), .Q(Q[0]), .QN(n117) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n44) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n136), .A2(n39), .B1(n47), .B2(n101), .ZN(n16) );
  INV_X1 U20 ( .A(D[19]), .ZN(n101) );
  OAI22_X1 U21 ( .A1(n129), .A2(n40), .B1(n45), .B2(n100), .ZN(n23) );
  INV_X1 U22 ( .A(D[12]), .ZN(n100) );
  OAI22_X1 U23 ( .A1(n130), .A2(n40), .B1(n45), .B2(n99), .ZN(n22) );
  INV_X1 U24 ( .A(D[13]), .ZN(n99) );
  OAI22_X1 U25 ( .A1(n131), .A2(n39), .B1(n46), .B2(n98), .ZN(n21) );
  INV_X1 U26 ( .A(D[14]), .ZN(n98) );
  OAI22_X1 U27 ( .A1(n132), .A2(n39), .B1(n46), .B2(n65), .ZN(n20) );
  INV_X1 U28 ( .A(D[15]), .ZN(n65) );
  OAI22_X1 U29 ( .A1(n137), .A2(n39), .B1(n47), .B2(n108), .ZN(n15) );
  INV_X1 U30 ( .A(D[20]), .ZN(n108) );
  OAI22_X1 U31 ( .A1(n138), .A2(n39), .B1(n47), .B2(n107), .ZN(n14) );
  INV_X1 U32 ( .A(D[21]), .ZN(n107) );
  OAI22_X1 U33 ( .A1(n139), .A2(n39), .B1(n48), .B2(n106), .ZN(n13) );
  INV_X1 U34 ( .A(D[22]), .ZN(n106) );
  OAI22_X1 U35 ( .A1(n140), .A2(n39), .B1(n48), .B2(n105), .ZN(n12) );
  INV_X1 U36 ( .A(D[23]), .ZN(n105) );
  OAI22_X1 U37 ( .A1(n141), .A2(n39), .B1(n48), .B2(n112), .ZN(n11) );
  INV_X1 U38 ( .A(D[24]), .ZN(n112) );
  OAI22_X1 U39 ( .A1(n142), .A2(n39), .B1(n48), .B2(n111), .ZN(n10) );
  INV_X1 U40 ( .A(D[25]), .ZN(n111) );
  OAI22_X1 U41 ( .A1(n143), .A2(n40), .B1(n41), .B2(n110), .ZN(n9) );
  INV_X1 U42 ( .A(D[26]), .ZN(n110) );
  OAI22_X1 U43 ( .A1(n144), .A2(n39), .B1(n41), .B2(n109), .ZN(n8) );
  INV_X1 U44 ( .A(D[27]), .ZN(n109) );
  OAI22_X1 U45 ( .A1(n145), .A2(n40), .B1(n41), .B2(n116), .ZN(n7) );
  INV_X1 U46 ( .A(D[28]), .ZN(n116) );
  OAI22_X1 U47 ( .A1(n146), .A2(n39), .B1(n41), .B2(n115), .ZN(n6) );
  INV_X1 U48 ( .A(D[29]), .ZN(n115) );
  OAI22_X1 U49 ( .A1(n147), .A2(n40), .B1(n42), .B2(n114), .ZN(n5) );
  INV_X1 U50 ( .A(D[30]), .ZN(n114) );
  OAI22_X1 U51 ( .A1(n148), .A2(n39), .B1(n42), .B2(n113), .ZN(n4) );
  INV_X1 U52 ( .A(D[31]), .ZN(n113) );
  OAI22_X1 U53 ( .A1(n133), .A2(n39), .B1(n46), .B2(n104), .ZN(n19) );
  INV_X1 U54 ( .A(D[16]), .ZN(n104) );
  OAI22_X1 U55 ( .A1(n134), .A2(n39), .B1(n46), .B2(n103), .ZN(n18) );
  INV_X1 U56 ( .A(D[17]), .ZN(n103) );
  OAI22_X1 U57 ( .A1(n135), .A2(n39), .B1(n47), .B2(n102), .ZN(n17) );
  INV_X1 U58 ( .A(D[18]), .ZN(n102) );
  OAI22_X1 U59 ( .A1(n117), .A2(n40), .B1(n42), .B2(n56), .ZN(n35) );
  INV_X1 U60 ( .A(D[0]), .ZN(n56) );
  OAI22_X1 U61 ( .A1(n125), .A2(n40), .B1(n44), .B2(n64), .ZN(n27) );
  INV_X1 U62 ( .A(D[8]), .ZN(n64) );
  OAI22_X1 U63 ( .A1(n126), .A2(n40), .B1(n44), .B2(n63), .ZN(n26) );
  INV_X1 U64 ( .A(D[9]), .ZN(n63) );
  OAI22_X1 U65 ( .A1(n127), .A2(n40), .B1(n45), .B2(n62), .ZN(n25) );
  INV_X1 U66 ( .A(D[10]), .ZN(n62) );
  OAI22_X1 U67 ( .A1(n121), .A2(n40), .B1(n43), .B2(n60), .ZN(n31) );
  INV_X1 U68 ( .A(D[4]), .ZN(n60) );
  OAI22_X1 U69 ( .A1(n122), .A2(n40), .B1(n43), .B2(n59), .ZN(n30) );
  INV_X1 U70 ( .A(D[5]), .ZN(n59) );
  OAI22_X1 U71 ( .A1(n123), .A2(n40), .B1(n44), .B2(n58), .ZN(n29) );
  INV_X1 U72 ( .A(D[6]), .ZN(n58) );
  OAI22_X1 U73 ( .A1(n128), .A2(n40), .B1(n45), .B2(n61), .ZN(n24) );
  INV_X1 U74 ( .A(D[11]), .ZN(n61) );
  OAI22_X1 U75 ( .A1(n124), .A2(n40), .B1(n44), .B2(n57), .ZN(n28) );
  INV_X1 U76 ( .A(D[7]), .ZN(n57) );
  OAI22_X1 U77 ( .A1(n118), .A2(n39), .B1(n42), .B2(n55), .ZN(n34) );
  INV_X1 U78 ( .A(D[1]), .ZN(n55) );
  OAI22_X1 U79 ( .A1(n119), .A2(n40), .B1(n43), .B2(n54), .ZN(n33) );
  INV_X1 U80 ( .A(D[2]), .ZN(n54) );
  OAI22_X1 U81 ( .A1(n120), .A2(n40), .B1(n43), .B2(n53), .ZN(n32) );
  INV_X1 U82 ( .A(D[3]), .ZN(n53) );
endmodule


module REG_GEN_NBIT32_5 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n50), .Q(Q[31]), .QN(n148) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n50), .Q(Q[30]), .QN(n147) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n50), .Q(Q[29]), .QN(n146) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n50), .Q(Q[28]), .QN(n145) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n50), .Q(Q[27]), .QN(n144) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n50), .Q(Q[26]), .QN(n143) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n50), .Q(Q[25]), .QN(n142) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n50), .Q(Q[24]), .QN(n141) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n50), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n50), .Q(Q[22]), .QN(n139) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n50), .Q(Q[21]), .QN(n138) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n50), .Q(Q[20]), .QN(n137) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n136) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n135) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n51), .Q(Q[17]), .QN(n134) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n133) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n132) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n131) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n51), .Q(Q[13]), .QN(n130) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n51), .Q(Q[12]), .QN(n129) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n51), .Q(Q[11]), .QN(n128) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n51), .Q(Q[10]), .QN(n127) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n51), .Q(Q[9]), .QN(n126) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n51), .Q(Q[8]), .QN(n125) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n52), .Q(Q[7]), .QN(n124) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n52), .Q(Q[6]), .QN(n123) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n52), .Q(Q[5]), .QN(n122) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n52), .Q(Q[4]), .QN(n121) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n52), .Q(Q[3]), .QN(n120) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n52), .Q(Q[2]), .QN(n119) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n52), .Q(Q[1]), .QN(n118) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n52), .Q(Q[0]), .QN(n117) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n44) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n117), .A2(n40), .B1(n42), .B2(n116), .ZN(n35) );
  INV_X1 U20 ( .A(D[0]), .ZN(n116) );
  OAI22_X1 U21 ( .A1(n118), .A2(n39), .B1(n42), .B2(n115), .ZN(n34) );
  INV_X1 U22 ( .A(D[1]), .ZN(n115) );
  OAI22_X1 U23 ( .A1(n143), .A2(n40), .B1(n41), .B2(n58), .ZN(n9) );
  INV_X1 U24 ( .A(D[26]), .ZN(n58) );
  OAI22_X1 U25 ( .A1(n144), .A2(n39), .B1(n41), .B2(n57), .ZN(n8) );
  INV_X1 U26 ( .A(D[27]), .ZN(n57) );
  OAI22_X1 U27 ( .A1(n145), .A2(n40), .B1(n41), .B2(n56), .ZN(n7) );
  INV_X1 U28 ( .A(D[28]), .ZN(n56) );
  OAI22_X1 U29 ( .A1(n146), .A2(n39), .B1(n41), .B2(n55), .ZN(n6) );
  INV_X1 U30 ( .A(D[29]), .ZN(n55) );
  OAI22_X1 U31 ( .A1(n147), .A2(n40), .B1(n42), .B2(n54), .ZN(n5) );
  INV_X1 U32 ( .A(D[30]), .ZN(n54) );
  OAI22_X1 U33 ( .A1(n148), .A2(n39), .B1(n42), .B2(n53), .ZN(n4) );
  INV_X1 U34 ( .A(D[31]), .ZN(n53) );
  OAI22_X1 U35 ( .A1(n119), .A2(n40), .B1(n43), .B2(n114), .ZN(n33) );
  INV_X1 U36 ( .A(D[2]), .ZN(n114) );
  OAI22_X1 U37 ( .A1(n120), .A2(n40), .B1(n43), .B2(n113), .ZN(n32) );
  INV_X1 U38 ( .A(D[3]), .ZN(n113) );
  OAI22_X1 U39 ( .A1(n121), .A2(n40), .B1(n43), .B2(n112), .ZN(n31) );
  INV_X1 U40 ( .A(D[4]), .ZN(n112) );
  OAI22_X1 U41 ( .A1(n122), .A2(n40), .B1(n43), .B2(n111), .ZN(n30) );
  INV_X1 U42 ( .A(D[5]), .ZN(n111) );
  OAI22_X1 U43 ( .A1(n123), .A2(n40), .B1(n44), .B2(n110), .ZN(n29) );
  INV_X1 U44 ( .A(D[6]), .ZN(n110) );
  OAI22_X1 U45 ( .A1(n124), .A2(n40), .B1(n44), .B2(n109), .ZN(n28) );
  INV_X1 U46 ( .A(D[7]), .ZN(n109) );
  OAI22_X1 U47 ( .A1(n125), .A2(n40), .B1(n44), .B2(n108), .ZN(n27) );
  INV_X1 U48 ( .A(D[8]), .ZN(n108) );
  OAI22_X1 U49 ( .A1(n126), .A2(n40), .B1(n44), .B2(n107), .ZN(n26) );
  INV_X1 U50 ( .A(D[9]), .ZN(n107) );
  OAI22_X1 U51 ( .A1(n127), .A2(n40), .B1(n45), .B2(n106), .ZN(n25) );
  INV_X1 U52 ( .A(D[10]), .ZN(n106) );
  OAI22_X1 U53 ( .A1(n128), .A2(n40), .B1(n45), .B2(n105), .ZN(n24) );
  INV_X1 U54 ( .A(D[11]), .ZN(n105) );
  OAI22_X1 U55 ( .A1(n129), .A2(n40), .B1(n45), .B2(n104), .ZN(n23) );
  INV_X1 U56 ( .A(D[12]), .ZN(n104) );
  OAI22_X1 U57 ( .A1(n130), .A2(n40), .B1(n45), .B2(n103), .ZN(n22) );
  INV_X1 U58 ( .A(D[13]), .ZN(n103) );
  OAI22_X1 U59 ( .A1(n131), .A2(n39), .B1(n46), .B2(n102), .ZN(n21) );
  INV_X1 U60 ( .A(D[14]), .ZN(n102) );
  OAI22_X1 U61 ( .A1(n132), .A2(n39), .B1(n46), .B2(n101), .ZN(n20) );
  INV_X1 U62 ( .A(D[15]), .ZN(n101) );
  OAI22_X1 U63 ( .A1(n133), .A2(n39), .B1(n46), .B2(n100), .ZN(n19) );
  INV_X1 U64 ( .A(D[16]), .ZN(n100) );
  OAI22_X1 U65 ( .A1(n134), .A2(n39), .B1(n46), .B2(n99), .ZN(n18) );
  INV_X1 U66 ( .A(D[17]), .ZN(n99) );
  OAI22_X1 U67 ( .A1(n135), .A2(n39), .B1(n47), .B2(n98), .ZN(n17) );
  INV_X1 U68 ( .A(D[18]), .ZN(n98) );
  OAI22_X1 U69 ( .A1(n136), .A2(n39), .B1(n47), .B2(n65), .ZN(n16) );
  INV_X1 U70 ( .A(D[19]), .ZN(n65) );
  OAI22_X1 U71 ( .A1(n137), .A2(n39), .B1(n47), .B2(n64), .ZN(n15) );
  INV_X1 U72 ( .A(D[20]), .ZN(n64) );
  OAI22_X1 U73 ( .A1(n138), .A2(n39), .B1(n47), .B2(n63), .ZN(n14) );
  INV_X1 U74 ( .A(D[21]), .ZN(n63) );
  OAI22_X1 U75 ( .A1(n139), .A2(n39), .B1(n48), .B2(n62), .ZN(n13) );
  INV_X1 U76 ( .A(D[22]), .ZN(n62) );
  OAI22_X1 U77 ( .A1(n140), .A2(n39), .B1(n48), .B2(n61), .ZN(n12) );
  INV_X1 U78 ( .A(D[23]), .ZN(n61) );
  OAI22_X1 U79 ( .A1(n141), .A2(n39), .B1(n48), .B2(n60), .ZN(n11) );
  INV_X1 U80 ( .A(D[24]), .ZN(n60) );
  OAI22_X1 U81 ( .A1(n142), .A2(n39), .B1(n48), .B2(n59), .ZN(n10) );
  INV_X1 U82 ( .A(D[25]), .ZN(n59) );
endmodule


module REG_GEN_NBIT32_4 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  DFFR_X1 \Q_reg[31]  ( .D(n4), .CK(CK), .RN(n52), .Q(Q[31]), .QN(n148) );
  DFFR_X1 \Q_reg[30]  ( .D(n5), .CK(CK), .RN(n52), .Q(Q[30]), .QN(n147) );
  DFFR_X1 \Q_reg[29]  ( .D(n6), .CK(CK), .RN(n52), .Q(Q[29]), .QN(n146) );
  DFFR_X1 \Q_reg[28]  ( .D(n7), .CK(CK), .RN(n52), .Q(Q[28]), .QN(n145) );
  DFFR_X1 \Q_reg[27]  ( .D(n8), .CK(CK), .RN(n52), .Q(Q[27]), .QN(n144) );
  DFFR_X1 \Q_reg[26]  ( .D(n9), .CK(CK), .RN(n52), .Q(Q[26]), .QN(n143) );
  DFFR_X1 \Q_reg[25]  ( .D(n10), .CK(CK), .RN(n52), .Q(Q[25]), .QN(n142) );
  DFFR_X1 \Q_reg[24]  ( .D(n11), .CK(CK), .RN(n52), .Q(Q[24]), .QN(n141) );
  DFFR_X1 \Q_reg[23]  ( .D(n12), .CK(CK), .RN(n51), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n13), .CK(CK), .RN(n51), .Q(Q[22]), .QN(n139) );
  DFFR_X1 \Q_reg[21]  ( .D(n14), .CK(CK), .RN(n51), .Q(Q[21]), .QN(n138) );
  DFFR_X1 \Q_reg[20]  ( .D(n15), .CK(CK), .RN(n51), .Q(Q[20]), .QN(n137) );
  DFFR_X1 \Q_reg[19]  ( .D(n16), .CK(CK), .RN(n51), .Q(Q[19]), .QN(n136) );
  DFFR_X1 \Q_reg[18]  ( .D(n17), .CK(CK), .RN(n51), .Q(Q[18]), .QN(n135) );
  DFFR_X1 \Q_reg[17]  ( .D(n18), .CK(CK), .RN(n51), .Q(Q[17]), .QN(n134) );
  DFFR_X1 \Q_reg[16]  ( .D(n19), .CK(CK), .RN(n51), .Q(Q[16]), .QN(n133) );
  DFFR_X1 \Q_reg[15]  ( .D(n20), .CK(CK), .RN(n51), .Q(Q[15]), .QN(n132) );
  DFFR_X1 \Q_reg[14]  ( .D(n21), .CK(CK), .RN(n51), .Q(Q[14]), .QN(n131) );
  DFFR_X1 \Q_reg[13]  ( .D(n22), .CK(CK), .RN(n51), .Q(Q[13]), .QN(n130) );
  DFFR_X1 \Q_reg[12]  ( .D(n23), .CK(CK), .RN(n51), .Q(Q[12]), .QN(n129) );
  DFFR_X1 \Q_reg[11]  ( .D(n24), .CK(CK), .RN(n50), .Q(Q[11]), .QN(n128) );
  DFFR_X1 \Q_reg[10]  ( .D(n25), .CK(CK), .RN(n50), .Q(Q[10]), .QN(n127) );
  DFFR_X1 \Q_reg[9]  ( .D(n26), .CK(CK), .RN(n50), .Q(Q[9]), .QN(n126) );
  DFFR_X1 \Q_reg[8]  ( .D(n27), .CK(CK), .RN(n50), .Q(Q[8]), .QN(n125) );
  DFFR_X1 \Q_reg[7]  ( .D(n28), .CK(CK), .RN(n50), .Q(Q[7]), .QN(n124) );
  DFFR_X1 \Q_reg[6]  ( .D(n29), .CK(CK), .RN(n50), .Q(Q[6]), .QN(n123) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CK), .RN(n50), .Q(Q[5]), .QN(n122) );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(CK), .RN(n50), .Q(Q[4]), .QN(n121) );
  DFFR_X1 \Q_reg[3]  ( .D(n32), .CK(CK), .RN(n50), .Q(Q[3]), .QN(n120) );
  DFFR_X1 \Q_reg[2]  ( .D(n33), .CK(CK), .RN(n50), .Q(Q[2]), .QN(n119) );
  DFFR_X1 \Q_reg[1]  ( .D(n34), .CK(CK), .RN(n50), .Q(Q[1]), .QN(n118) );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(CK), .RN(n50), .Q(Q[0]), .QN(n117) );
  INV_X1 U2 ( .A(n49), .ZN(n40) );
  INV_X1 U3 ( .A(n49), .ZN(n39) );
  BUF_X1 U4 ( .A(RESET_n), .Z(n50) );
  BUF_X1 U5 ( .A(RESET_n), .Z(n51) );
  BUF_X1 U6 ( .A(RESET_n), .Z(n52) );
  BUF_X1 U7 ( .A(n38), .Z(n49) );
  BUF_X1 U8 ( .A(n36), .Z(n43) );
  BUF_X1 U9 ( .A(n37), .Z(n44) );
  BUF_X1 U10 ( .A(n37), .Z(n45) );
  BUF_X1 U11 ( .A(n37), .Z(n46) );
  BUF_X1 U12 ( .A(n38), .Z(n47) );
  BUF_X1 U13 ( .A(n38), .Z(n48) );
  BUF_X1 U14 ( .A(n36), .Z(n41) );
  BUF_X1 U15 ( .A(n36), .Z(n42) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n38) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n37) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n36) );
  OAI22_X1 U19 ( .A1(n117), .A2(n40), .B1(n42), .B2(n116), .ZN(n35) );
  INV_X1 U20 ( .A(D[0]), .ZN(n116) );
  OAI22_X1 U21 ( .A1(n118), .A2(n39), .B1(n42), .B2(n115), .ZN(n34) );
  INV_X1 U22 ( .A(D[1]), .ZN(n115) );
  OAI22_X1 U23 ( .A1(n143), .A2(n40), .B1(n41), .B2(n58), .ZN(n9) );
  INV_X1 U24 ( .A(D[26]), .ZN(n58) );
  OAI22_X1 U25 ( .A1(n144), .A2(n39), .B1(n41), .B2(n57), .ZN(n8) );
  INV_X1 U26 ( .A(D[27]), .ZN(n57) );
  OAI22_X1 U27 ( .A1(n145), .A2(n40), .B1(n41), .B2(n56), .ZN(n7) );
  INV_X1 U28 ( .A(D[28]), .ZN(n56) );
  OAI22_X1 U29 ( .A1(n146), .A2(n39), .B1(n41), .B2(n55), .ZN(n6) );
  INV_X1 U30 ( .A(D[29]), .ZN(n55) );
  OAI22_X1 U31 ( .A1(n147), .A2(n40), .B1(n42), .B2(n54), .ZN(n5) );
  INV_X1 U32 ( .A(D[30]), .ZN(n54) );
  OAI22_X1 U33 ( .A1(n148), .A2(n39), .B1(n42), .B2(n53), .ZN(n4) );
  INV_X1 U34 ( .A(D[31]), .ZN(n53) );
  OAI22_X1 U35 ( .A1(n129), .A2(n40), .B1(n45), .B2(n104), .ZN(n23) );
  INV_X1 U36 ( .A(D[12]), .ZN(n104) );
  OAI22_X1 U37 ( .A1(n130), .A2(n40), .B1(n45), .B2(n103), .ZN(n22) );
  INV_X1 U38 ( .A(D[13]), .ZN(n103) );
  OAI22_X1 U39 ( .A1(n131), .A2(n39), .B1(n46), .B2(n102), .ZN(n21) );
  INV_X1 U40 ( .A(D[14]), .ZN(n102) );
  OAI22_X1 U41 ( .A1(n132), .A2(n39), .B1(n46), .B2(n101), .ZN(n20) );
  INV_X1 U42 ( .A(D[15]), .ZN(n101) );
  OAI22_X1 U43 ( .A1(n133), .A2(n39), .B1(n46), .B2(n100), .ZN(n19) );
  INV_X1 U44 ( .A(D[16]), .ZN(n100) );
  OAI22_X1 U45 ( .A1(n134), .A2(n39), .B1(n46), .B2(n99), .ZN(n18) );
  INV_X1 U46 ( .A(D[17]), .ZN(n99) );
  OAI22_X1 U47 ( .A1(n135), .A2(n39), .B1(n47), .B2(n98), .ZN(n17) );
  INV_X1 U48 ( .A(D[18]), .ZN(n98) );
  OAI22_X1 U49 ( .A1(n136), .A2(n39), .B1(n47), .B2(n65), .ZN(n16) );
  INV_X1 U50 ( .A(D[19]), .ZN(n65) );
  OAI22_X1 U51 ( .A1(n137), .A2(n39), .B1(n47), .B2(n64), .ZN(n15) );
  INV_X1 U52 ( .A(D[20]), .ZN(n64) );
  OAI22_X1 U53 ( .A1(n138), .A2(n39), .B1(n47), .B2(n63), .ZN(n14) );
  INV_X1 U54 ( .A(D[21]), .ZN(n63) );
  OAI22_X1 U55 ( .A1(n139), .A2(n39), .B1(n48), .B2(n62), .ZN(n13) );
  INV_X1 U56 ( .A(D[22]), .ZN(n62) );
  OAI22_X1 U57 ( .A1(n140), .A2(n39), .B1(n48), .B2(n61), .ZN(n12) );
  INV_X1 U58 ( .A(D[23]), .ZN(n61) );
  OAI22_X1 U59 ( .A1(n141), .A2(n39), .B1(n48), .B2(n60), .ZN(n11) );
  INV_X1 U60 ( .A(D[24]), .ZN(n60) );
  OAI22_X1 U61 ( .A1(n142), .A2(n39), .B1(n48), .B2(n59), .ZN(n10) );
  INV_X1 U62 ( .A(D[25]), .ZN(n59) );
  OAI22_X1 U63 ( .A1(n119), .A2(n40), .B1(n43), .B2(n114), .ZN(n33) );
  INV_X1 U64 ( .A(D[2]), .ZN(n114) );
  OAI22_X1 U65 ( .A1(n120), .A2(n40), .B1(n43), .B2(n113), .ZN(n32) );
  INV_X1 U66 ( .A(D[3]), .ZN(n113) );
  OAI22_X1 U67 ( .A1(n121), .A2(n40), .B1(n43), .B2(n112), .ZN(n31) );
  INV_X1 U68 ( .A(D[4]), .ZN(n112) );
  OAI22_X1 U69 ( .A1(n122), .A2(n40), .B1(n43), .B2(n111), .ZN(n30) );
  INV_X1 U70 ( .A(D[5]), .ZN(n111) );
  OAI22_X1 U71 ( .A1(n123), .A2(n40), .B1(n44), .B2(n110), .ZN(n29) );
  INV_X1 U72 ( .A(D[6]), .ZN(n110) );
  OAI22_X1 U73 ( .A1(n124), .A2(n40), .B1(n44), .B2(n109), .ZN(n28) );
  INV_X1 U74 ( .A(D[7]), .ZN(n109) );
  OAI22_X1 U75 ( .A1(n125), .A2(n40), .B1(n44), .B2(n108), .ZN(n27) );
  INV_X1 U76 ( .A(D[8]), .ZN(n108) );
  OAI22_X1 U77 ( .A1(n126), .A2(n40), .B1(n44), .B2(n107), .ZN(n26) );
  INV_X1 U78 ( .A(D[9]), .ZN(n107) );
  OAI22_X1 U79 ( .A1(n127), .A2(n40), .B1(n45), .B2(n106), .ZN(n25) );
  INV_X1 U80 ( .A(D[10]), .ZN(n106) );
  OAI22_X1 U81 ( .A1(n128), .A2(n40), .B1(n45), .B2(n105), .ZN(n24) );
  INV_X1 U82 ( .A(D[11]), .ZN(n105) );
endmodule


module executionUnit_nbit32 ( r1, r2, imm, j_lab, pc, RW_R, RW_I, s2, s3, rst, 
        clk, en_reg, alu_sel, alu_out, alu_fw_out, r2_out, b_lab_out, 
        pc_exe_out, rw_exe, j_lab_out );
  input [31:0] r1;
  input [31:0] r2;
  input [31:0] imm;
  input [31:0] j_lab;
  input [31:0] pc;
  input [31:0] RW_R;
  input [31:0] RW_I;
  input [3:0] alu_sel;
  output [31:0] alu_out;
  output [31:0] alu_fw_out;
  output [31:0] r2_out;
  output [31:0] b_lab_out;
  output [31:0] pc_exe_out;
  output [31:0] rw_exe;
  output [31:0] j_lab_out;
  input s2, s3, rst, clk, en_reg;
  wire   n1, n2;
  wire   [31:0] mux_out;
  wire   [31:0] rw_s;
  wire   [31:0] pc_b;
  wire   [31:0] pc_j;

  MUX21_GENERIC_NBIT32_8 lo_mux ( .A(r2), .B(imm), .SEL(s2), .Y(mux_out) );
  MUX21_GENERIC_NBIT32_7 RW_mux ( .A(RW_R), .B(RW_I), .SEL(s3), .Y(rw_s) );
  alu alu_dut ( .data_in1({r1[31:26], n1, r1[24:0]}), .data_in2(mux_out), 
        .op_sel(alu_sel), .data_out(alu_fw_out) );
  REG_GEN_NBIT32_9 reg_alu ( .D(alu_fw_out), .CK(clk), .Enable_n(n2), 
        .RESET_n(rst), .Q(alu_out) );
  REG_GEN_NBIT32_8 ls_reg ( .D(r2), .CK(clk), .Enable_n(n2), .RESET_n(rst), 
        .Q(r2_out) );
  P4_ADDER_NBIT32_NBIT_PER_BLOCK4_3 pc_br ( .A(imm), .B(pc), .Cin(1'b0), .Y(
        pc_b) );
  P4_ADDER_NBIT32_NBIT_PER_BLOCK4_2 pc_jp ( .A(j_lab), .B(pc), .Cin(1'b0), .Y(
        pc_j) );
  REG_GEN_NBIT32_7 pc_reg_b ( .D(pc_b), .CK(clk), .Enable_n(n2), .RESET_n(rst), 
        .Q(b_lab_out) );
  REG_GEN_NBIT32_6 pc_reg_j ( .D(pc_j), .CK(clk), .Enable_n(n2), .RESET_n(rst), 
        .Q(j_lab_out) );
  REG_GEN_NBIT32_5 pc_reg ( .D(pc), .CK(clk), .Enable_n(n2), .RESET_n(rst), 
        .Q(pc_exe_out) );
  REG_GEN_NBIT32_4 rw_reg ( .D(rw_s), .CK(clk), .Enable_n(n2), .RESET_n(rst), 
        .Q(rw_exe) );
  BUF_X1 U2 ( .A(r1[25]), .Z(n1) );
  BUF_X1 U3 ( .A(en_reg), .Z(n2) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n33, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142;

  INV_X1 U1 ( .A(n78), .ZN(n68) );
  INV_X1 U2 ( .A(n78), .ZN(n69) );
  BUF_X1 U3 ( .A(n33), .Z(n70) );
  BUF_X1 U4 ( .A(n67), .Z(n76) );
  BUF_X1 U5 ( .A(n66), .Z(n75) );
  BUF_X1 U6 ( .A(n66), .Z(n73) );
  BUF_X1 U7 ( .A(n33), .Z(n72) );
  BUF_X1 U8 ( .A(n66), .Z(n74) );
  BUF_X1 U9 ( .A(n33), .Z(n71) );
  BUF_X1 U10 ( .A(n67), .Z(n78) );
  BUF_X1 U11 ( .A(n67), .Z(n77) );
  BUF_X1 U12 ( .A(SEL), .Z(n67) );
  BUF_X1 U13 ( .A(SEL), .Z(n66) );
  BUF_X1 U14 ( .A(SEL), .Z(n33) );
  INV_X1 U15 ( .A(n142), .ZN(Y[9]) );
  AOI22_X1 U16 ( .A1(A[9]), .A2(n68), .B1(n77), .B2(B[9]), .ZN(n142) );
  INV_X1 U17 ( .A(n111), .ZN(Y[0]) );
  AOI22_X1 U18 ( .A1(A[0]), .A2(n68), .B1(B[0]), .B2(n77), .ZN(n111) );
  INV_X1 U19 ( .A(n122), .ZN(Y[1]) );
  AOI22_X1 U20 ( .A1(A[1]), .A2(n68), .B1(B[1]), .B2(n74), .ZN(n122) );
  INV_X1 U21 ( .A(n133), .ZN(Y[2]) );
  AOI22_X1 U22 ( .A1(A[2]), .A2(n69), .B1(B[2]), .B2(n71), .ZN(n133) );
  INV_X1 U23 ( .A(n136), .ZN(Y[3]) );
  AOI22_X1 U24 ( .A1(A[3]), .A2(n69), .B1(B[3]), .B2(n71), .ZN(n136) );
  INV_X1 U25 ( .A(n137), .ZN(Y[4]) );
  AOI22_X1 U26 ( .A1(A[4]), .A2(n68), .B1(B[4]), .B2(n71), .ZN(n137) );
  INV_X1 U27 ( .A(n138), .ZN(Y[5]) );
  AOI22_X1 U28 ( .A1(A[5]), .A2(n69), .B1(B[5]), .B2(n70), .ZN(n138) );
  INV_X1 U29 ( .A(n139), .ZN(Y[6]) );
  AOI22_X1 U30 ( .A1(A[6]), .A2(n68), .B1(B[6]), .B2(n70), .ZN(n139) );
  INV_X1 U31 ( .A(n140), .ZN(Y[7]) );
  AOI22_X1 U32 ( .A1(A[7]), .A2(n69), .B1(B[7]), .B2(n70), .ZN(n140) );
  INV_X1 U33 ( .A(n141), .ZN(Y[8]) );
  AOI22_X1 U34 ( .A1(A[8]), .A2(n68), .B1(B[8]), .B2(n70), .ZN(n141) );
  INV_X1 U35 ( .A(n112), .ZN(Y[10]) );
  AOI22_X1 U36 ( .A1(A[10]), .A2(n68), .B1(B[10]), .B2(n77), .ZN(n112) );
  INV_X1 U37 ( .A(n113), .ZN(Y[11]) );
  AOI22_X1 U38 ( .A1(A[11]), .A2(n68), .B1(B[11]), .B2(n77), .ZN(n113) );
  INV_X1 U39 ( .A(n114), .ZN(Y[12]) );
  AOI22_X1 U40 ( .A1(A[12]), .A2(n68), .B1(B[12]), .B2(n76), .ZN(n114) );
  INV_X1 U41 ( .A(n115), .ZN(Y[13]) );
  AOI22_X1 U42 ( .A1(A[13]), .A2(n68), .B1(B[13]), .B2(n76), .ZN(n115) );
  INV_X1 U43 ( .A(n116), .ZN(Y[14]) );
  AOI22_X1 U44 ( .A1(A[14]), .A2(n68), .B1(B[14]), .B2(n76), .ZN(n116) );
  INV_X1 U45 ( .A(n117), .ZN(Y[15]) );
  AOI22_X1 U46 ( .A1(A[15]), .A2(n68), .B1(B[15]), .B2(n76), .ZN(n117) );
  INV_X1 U47 ( .A(n118), .ZN(Y[16]) );
  AOI22_X1 U48 ( .A1(A[16]), .A2(n68), .B1(B[16]), .B2(n75), .ZN(n118) );
  INV_X1 U49 ( .A(n119), .ZN(Y[17]) );
  AOI22_X1 U50 ( .A1(A[17]), .A2(n68), .B1(B[17]), .B2(n75), .ZN(n119) );
  INV_X1 U51 ( .A(n120), .ZN(Y[18]) );
  AOI22_X1 U52 ( .A1(A[18]), .A2(n68), .B1(B[18]), .B2(n75), .ZN(n120) );
  INV_X1 U53 ( .A(n121), .ZN(Y[19]) );
  AOI22_X1 U54 ( .A1(A[19]), .A2(n68), .B1(B[19]), .B2(n75), .ZN(n121) );
  INV_X1 U55 ( .A(n123), .ZN(Y[20]) );
  AOI22_X1 U56 ( .A1(A[20]), .A2(n69), .B1(B[20]), .B2(n74), .ZN(n123) );
  INV_X1 U57 ( .A(n124), .ZN(Y[21]) );
  AOI22_X1 U58 ( .A1(A[21]), .A2(n69), .B1(B[21]), .B2(n74), .ZN(n124) );
  INV_X1 U59 ( .A(n125), .ZN(Y[22]) );
  AOI22_X1 U60 ( .A1(A[22]), .A2(n69), .B1(B[22]), .B2(n73), .ZN(n125) );
  INV_X1 U61 ( .A(n126), .ZN(Y[23]) );
  AOI22_X1 U62 ( .A1(A[23]), .A2(n69), .B1(B[23]), .B2(n73), .ZN(n126) );
  INV_X1 U63 ( .A(n127), .ZN(Y[24]) );
  AOI22_X1 U64 ( .A1(A[24]), .A2(n69), .B1(B[24]), .B2(n73), .ZN(n127) );
  INV_X1 U65 ( .A(n128), .ZN(Y[25]) );
  AOI22_X1 U66 ( .A1(A[25]), .A2(n69), .B1(B[25]), .B2(n73), .ZN(n128) );
  INV_X1 U67 ( .A(n129), .ZN(Y[26]) );
  AOI22_X1 U68 ( .A1(A[26]), .A2(n69), .B1(B[26]), .B2(n72), .ZN(n129) );
  INV_X1 U69 ( .A(n130), .ZN(Y[27]) );
  AOI22_X1 U70 ( .A1(A[27]), .A2(n69), .B1(B[27]), .B2(n72), .ZN(n130) );
  INV_X1 U71 ( .A(n131), .ZN(Y[28]) );
  AOI22_X1 U72 ( .A1(A[28]), .A2(n69), .B1(B[28]), .B2(n72), .ZN(n131) );
  INV_X1 U73 ( .A(n132), .ZN(Y[29]) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n69), .B1(B[29]), .B2(n72), .ZN(n132) );
  INV_X1 U75 ( .A(n134), .ZN(Y[30]) );
  AOI22_X1 U76 ( .A1(A[30]), .A2(n69), .B1(B[30]), .B2(n74), .ZN(n134) );
  INV_X1 U77 ( .A(n135), .ZN(Y[31]) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n69), .B1(B[31]), .B2(n71), .ZN(n135) );
endmodule


module branch_block_nbit32 ( branch_op, cmp_out, PC, label_PC, next_PC );
  input [31:0] cmp_out;
  input [31:0] PC;
  input [31:0] label_PC;
  output [31:0] next_PC;
  input branch_op;
  wire   branch_taken;

  MUX21_GENERIC_NBIT32_1 next_pc_mux ( .A(PC), .B(label_PC), .SEL(branch_taken), .Y(next_PC) );
  AND2_X1 U1 ( .A1(cmp_out[0]), .A2(branch_op), .ZN(branch_taken) );
endmodule


module MUX21_GENERIC_NBIT32_6 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n33, n66, n67, n100;

  BUF_X1 U1 ( .A(n100), .Z(n33) );
  BUF_X1 U2 ( .A(n100), .Z(n66) );
  BUF_X1 U3 ( .A(n100), .Z(n67) );
  INV_X1 U4 ( .A(n34), .ZN(Y[9]) );
  AOI22_X1 U5 ( .A1(A[9]), .A2(n67), .B1(SEL), .B2(B[9]), .ZN(n34) );
  INV_X1 U6 ( .A(n65), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(n33), .B1(B[0]), .B2(SEL), .ZN(n65) );
  INV_X1 U8 ( .A(n54), .ZN(Y[1]) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n33), .B1(B[1]), .B2(SEL), .ZN(n54) );
  INV_X1 U10 ( .A(n43), .ZN(Y[2]) );
  AOI22_X1 U11 ( .A1(A[2]), .A2(n66), .B1(B[2]), .B2(SEL), .ZN(n43) );
  INV_X1 U12 ( .A(n40), .ZN(Y[3]) );
  AOI22_X1 U13 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(SEL), .ZN(n40) );
  INV_X1 U14 ( .A(n39), .ZN(Y[4]) );
  AOI22_X1 U15 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(SEL), .ZN(n39) );
  INV_X1 U16 ( .A(n38), .ZN(Y[5]) );
  AOI22_X1 U17 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(SEL), .ZN(n38) );
  INV_X1 U18 ( .A(n37), .ZN(Y[6]) );
  AOI22_X1 U19 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(SEL), .ZN(n37) );
  INV_X1 U20 ( .A(n36), .ZN(Y[7]) );
  AOI22_X1 U21 ( .A1(A[7]), .A2(n67), .B1(B[7]), .B2(SEL), .ZN(n36) );
  INV_X1 U22 ( .A(n35), .ZN(Y[8]) );
  AOI22_X1 U23 ( .A1(A[8]), .A2(n67), .B1(B[8]), .B2(SEL), .ZN(n35) );
  INV_X1 U24 ( .A(n64), .ZN(Y[10]) );
  AOI22_X1 U25 ( .A1(A[10]), .A2(n33), .B1(B[10]), .B2(SEL), .ZN(n64) );
  INV_X1 U26 ( .A(n63), .ZN(Y[11]) );
  AOI22_X1 U27 ( .A1(A[11]), .A2(n33), .B1(B[11]), .B2(SEL), .ZN(n63) );
  INV_X1 U28 ( .A(n62), .ZN(Y[12]) );
  AOI22_X1 U29 ( .A1(A[12]), .A2(n33), .B1(B[12]), .B2(SEL), .ZN(n62) );
  INV_X1 U30 ( .A(n61), .ZN(Y[13]) );
  AOI22_X1 U31 ( .A1(A[13]), .A2(n33), .B1(B[13]), .B2(SEL), .ZN(n61) );
  INV_X1 U32 ( .A(n60), .ZN(Y[14]) );
  AOI22_X1 U33 ( .A1(A[14]), .A2(n33), .B1(B[14]), .B2(SEL), .ZN(n60) );
  INV_X1 U34 ( .A(n59), .ZN(Y[15]) );
  AOI22_X1 U35 ( .A1(A[15]), .A2(n33), .B1(B[15]), .B2(SEL), .ZN(n59) );
  INV_X1 U36 ( .A(n58), .ZN(Y[16]) );
  AOI22_X1 U37 ( .A1(A[16]), .A2(n33), .B1(B[16]), .B2(SEL), .ZN(n58) );
  INV_X1 U38 ( .A(n57), .ZN(Y[17]) );
  AOI22_X1 U39 ( .A1(A[17]), .A2(n33), .B1(B[17]), .B2(SEL), .ZN(n57) );
  INV_X1 U40 ( .A(n56), .ZN(Y[18]) );
  AOI22_X1 U41 ( .A1(A[18]), .A2(n33), .B1(B[18]), .B2(SEL), .ZN(n56) );
  INV_X1 U42 ( .A(n55), .ZN(Y[19]) );
  AOI22_X1 U43 ( .A1(A[19]), .A2(n33), .B1(B[19]), .B2(SEL), .ZN(n55) );
  INV_X1 U44 ( .A(n53), .ZN(Y[20]) );
  AOI22_X1 U45 ( .A1(A[20]), .A2(n66), .B1(B[20]), .B2(SEL), .ZN(n53) );
  INV_X1 U46 ( .A(n52), .ZN(Y[21]) );
  AOI22_X1 U47 ( .A1(A[21]), .A2(n66), .B1(B[21]), .B2(SEL), .ZN(n52) );
  INV_X1 U48 ( .A(n51), .ZN(Y[22]) );
  AOI22_X1 U49 ( .A1(A[22]), .A2(n66), .B1(B[22]), .B2(SEL), .ZN(n51) );
  INV_X1 U50 ( .A(n50), .ZN(Y[23]) );
  AOI22_X1 U51 ( .A1(A[23]), .A2(n66), .B1(B[23]), .B2(SEL), .ZN(n50) );
  INV_X1 U52 ( .A(n49), .ZN(Y[24]) );
  AOI22_X1 U53 ( .A1(A[24]), .A2(n66), .B1(B[24]), .B2(SEL), .ZN(n49) );
  INV_X1 U54 ( .A(n48), .ZN(Y[25]) );
  AOI22_X1 U55 ( .A1(A[25]), .A2(n66), .B1(B[25]), .B2(SEL), .ZN(n48) );
  INV_X1 U56 ( .A(n47), .ZN(Y[26]) );
  AOI22_X1 U57 ( .A1(A[26]), .A2(n66), .B1(B[26]), .B2(SEL), .ZN(n47) );
  INV_X1 U58 ( .A(n46), .ZN(Y[27]) );
  AOI22_X1 U59 ( .A1(A[27]), .A2(n66), .B1(B[27]), .B2(SEL), .ZN(n46) );
  INV_X1 U60 ( .A(n45), .ZN(Y[28]) );
  AOI22_X1 U61 ( .A1(A[28]), .A2(n66), .B1(B[28]), .B2(SEL), .ZN(n45) );
  INV_X1 U62 ( .A(n44), .ZN(Y[29]) );
  AOI22_X1 U63 ( .A1(A[29]), .A2(n66), .B1(B[29]), .B2(SEL), .ZN(n44) );
  INV_X1 U64 ( .A(n42), .ZN(Y[30]) );
  AOI22_X1 U65 ( .A1(A[30]), .A2(n66), .B1(B[30]), .B2(SEL), .ZN(n42) );
  INV_X1 U66 ( .A(n41), .ZN(Y[31]) );
  AOI22_X1 U67 ( .A1(A[31]), .A2(n67), .B1(B[31]), .B2(SEL), .ZN(n41) );
  INV_X1 U68 ( .A(SEL), .ZN(n100) );
endmodule


module MUX21_GENERIC_NBIT32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n33, n66, n67, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132;

  BUF_X1 U1 ( .A(n100), .Z(n33) );
  BUF_X1 U2 ( .A(n100), .Z(n66) );
  BUF_X1 U3 ( .A(n100), .Z(n67) );
  INV_X1 U4 ( .A(n101), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n33), .B1(B[0]), .B2(SEL), .ZN(n101) );
  INV_X1 U6 ( .A(n112), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n33), .B1(B[1]), .B2(SEL), .ZN(n112) );
  INV_X1 U8 ( .A(n116), .ZN(Y[23]) );
  AOI22_X1 U9 ( .A1(A[23]), .A2(n66), .B1(B[23]), .B2(SEL), .ZN(n116) );
  INV_X1 U10 ( .A(n117), .ZN(Y[24]) );
  AOI22_X1 U11 ( .A1(A[24]), .A2(n66), .B1(B[24]), .B2(SEL), .ZN(n117) );
  INV_X1 U12 ( .A(n118), .ZN(Y[25]) );
  AOI22_X1 U13 ( .A1(A[25]), .A2(n66), .B1(B[25]), .B2(SEL), .ZN(n118) );
  INV_X1 U14 ( .A(n119), .ZN(Y[26]) );
  AOI22_X1 U15 ( .A1(A[26]), .A2(n66), .B1(B[26]), .B2(SEL), .ZN(n119) );
  INV_X1 U16 ( .A(n120), .ZN(Y[27]) );
  AOI22_X1 U17 ( .A1(A[27]), .A2(n66), .B1(B[27]), .B2(SEL), .ZN(n120) );
  INV_X1 U18 ( .A(n121), .ZN(Y[28]) );
  AOI22_X1 U19 ( .A1(A[28]), .A2(n66), .B1(B[28]), .B2(SEL), .ZN(n121) );
  INV_X1 U20 ( .A(n123), .ZN(Y[2]) );
  AOI22_X1 U21 ( .A1(A[2]), .A2(n66), .B1(B[2]), .B2(SEL), .ZN(n123) );
  INV_X1 U22 ( .A(n126), .ZN(Y[3]) );
  AOI22_X1 U23 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(SEL), .ZN(n126) );
  INV_X1 U24 ( .A(n127), .ZN(Y[4]) );
  AOI22_X1 U25 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(SEL), .ZN(n127) );
  INV_X1 U26 ( .A(n128), .ZN(Y[5]) );
  AOI22_X1 U27 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(SEL), .ZN(n128) );
  INV_X1 U28 ( .A(n129), .ZN(Y[6]) );
  AOI22_X1 U29 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(SEL), .ZN(n129) );
  INV_X1 U30 ( .A(n130), .ZN(Y[7]) );
  AOI22_X1 U31 ( .A1(A[7]), .A2(n67), .B1(B[7]), .B2(SEL), .ZN(n130) );
  INV_X1 U32 ( .A(n131), .ZN(Y[8]) );
  AOI22_X1 U33 ( .A1(A[8]), .A2(n67), .B1(B[8]), .B2(SEL), .ZN(n131) );
  INV_X1 U34 ( .A(n132), .ZN(Y[9]) );
  AOI22_X1 U35 ( .A1(A[9]), .A2(n67), .B1(SEL), .B2(B[9]), .ZN(n132) );
  INV_X1 U36 ( .A(n102), .ZN(Y[10]) );
  AOI22_X1 U37 ( .A1(A[10]), .A2(n33), .B1(B[10]), .B2(SEL), .ZN(n102) );
  INV_X1 U38 ( .A(n103), .ZN(Y[11]) );
  AOI22_X1 U39 ( .A1(A[11]), .A2(n33), .B1(B[11]), .B2(SEL), .ZN(n103) );
  INV_X1 U40 ( .A(n104), .ZN(Y[12]) );
  AOI22_X1 U41 ( .A1(A[12]), .A2(n33), .B1(B[12]), .B2(SEL), .ZN(n104) );
  INV_X1 U42 ( .A(n105), .ZN(Y[13]) );
  AOI22_X1 U43 ( .A1(A[13]), .A2(n33), .B1(B[13]), .B2(SEL), .ZN(n105) );
  INV_X1 U44 ( .A(n106), .ZN(Y[14]) );
  AOI22_X1 U45 ( .A1(A[14]), .A2(n33), .B1(B[14]), .B2(SEL), .ZN(n106) );
  INV_X1 U46 ( .A(n107), .ZN(Y[15]) );
  AOI22_X1 U47 ( .A1(A[15]), .A2(n33), .B1(B[15]), .B2(SEL), .ZN(n107) );
  INV_X1 U48 ( .A(n108), .ZN(Y[16]) );
  AOI22_X1 U49 ( .A1(A[16]), .A2(n33), .B1(B[16]), .B2(SEL), .ZN(n108) );
  INV_X1 U50 ( .A(n109), .ZN(Y[17]) );
  AOI22_X1 U51 ( .A1(A[17]), .A2(n33), .B1(B[17]), .B2(SEL), .ZN(n109) );
  INV_X1 U52 ( .A(n110), .ZN(Y[18]) );
  AOI22_X1 U53 ( .A1(A[18]), .A2(n33), .B1(B[18]), .B2(SEL), .ZN(n110) );
  INV_X1 U54 ( .A(n111), .ZN(Y[19]) );
  AOI22_X1 U55 ( .A1(A[19]), .A2(n33), .B1(B[19]), .B2(SEL), .ZN(n111) );
  INV_X1 U56 ( .A(n113), .ZN(Y[20]) );
  AOI22_X1 U57 ( .A1(A[20]), .A2(n66), .B1(B[20]), .B2(SEL), .ZN(n113) );
  INV_X1 U58 ( .A(n114), .ZN(Y[21]) );
  AOI22_X1 U59 ( .A1(A[21]), .A2(n66), .B1(B[21]), .B2(SEL), .ZN(n114) );
  INV_X1 U60 ( .A(n115), .ZN(Y[22]) );
  AOI22_X1 U61 ( .A1(A[22]), .A2(n66), .B1(B[22]), .B2(SEL), .ZN(n115) );
  INV_X1 U62 ( .A(n122), .ZN(Y[29]) );
  AOI22_X1 U63 ( .A1(A[29]), .A2(n66), .B1(B[29]), .B2(SEL), .ZN(n122) );
  INV_X1 U64 ( .A(n124), .ZN(Y[30]) );
  AOI22_X1 U65 ( .A1(A[30]), .A2(n66), .B1(B[30]), .B2(SEL), .ZN(n124) );
  INV_X1 U66 ( .A(n125), .ZN(Y[31]) );
  AOI22_X1 U67 ( .A1(A[31]), .A2(n67), .B1(B[31]), .B2(SEL), .ZN(n125) );
  INV_X1 U68 ( .A(SEL), .ZN(n100) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n33, n66, n67, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132;

  BUF_X1 U1 ( .A(n100), .Z(n33) );
  BUF_X1 U2 ( .A(n100), .Z(n66) );
  BUF_X1 U3 ( .A(n100), .Z(n67) );
  INV_X1 U4 ( .A(n101), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n33), .B1(B[0]), .B2(SEL), .ZN(n101) );
  INV_X1 U6 ( .A(n112), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n33), .B1(B[1]), .B2(SEL), .ZN(n112) );
  INV_X1 U8 ( .A(n116), .ZN(Y[23]) );
  AOI22_X1 U9 ( .A1(A[23]), .A2(n66), .B1(B[23]), .B2(SEL), .ZN(n116) );
  INV_X1 U10 ( .A(n117), .ZN(Y[24]) );
  AOI22_X1 U11 ( .A1(A[24]), .A2(n66), .B1(B[24]), .B2(SEL), .ZN(n117) );
  INV_X1 U12 ( .A(n118), .ZN(Y[25]) );
  AOI22_X1 U13 ( .A1(A[25]), .A2(n66), .B1(B[25]), .B2(SEL), .ZN(n118) );
  INV_X1 U14 ( .A(n119), .ZN(Y[26]) );
  AOI22_X1 U15 ( .A1(A[26]), .A2(n66), .B1(B[26]), .B2(SEL), .ZN(n119) );
  INV_X1 U16 ( .A(n120), .ZN(Y[27]) );
  AOI22_X1 U17 ( .A1(A[27]), .A2(n66), .B1(B[27]), .B2(SEL), .ZN(n120) );
  INV_X1 U18 ( .A(n121), .ZN(Y[28]) );
  AOI22_X1 U19 ( .A1(A[28]), .A2(n66), .B1(B[28]), .B2(SEL), .ZN(n121) );
  INV_X1 U20 ( .A(n123), .ZN(Y[2]) );
  AOI22_X1 U21 ( .A1(A[2]), .A2(n66), .B1(B[2]), .B2(SEL), .ZN(n123) );
  INV_X1 U22 ( .A(n126), .ZN(Y[3]) );
  AOI22_X1 U23 ( .A1(A[3]), .A2(n67), .B1(B[3]), .B2(SEL), .ZN(n126) );
  INV_X1 U24 ( .A(n127), .ZN(Y[4]) );
  AOI22_X1 U25 ( .A1(A[4]), .A2(n67), .B1(B[4]), .B2(SEL), .ZN(n127) );
  INV_X1 U26 ( .A(n128), .ZN(Y[5]) );
  AOI22_X1 U27 ( .A1(A[5]), .A2(n67), .B1(B[5]), .B2(SEL), .ZN(n128) );
  INV_X1 U28 ( .A(n129), .ZN(Y[6]) );
  AOI22_X1 U29 ( .A1(A[6]), .A2(n67), .B1(B[6]), .B2(SEL), .ZN(n129) );
  INV_X1 U30 ( .A(n130), .ZN(Y[7]) );
  AOI22_X1 U31 ( .A1(A[7]), .A2(n67), .B1(B[7]), .B2(SEL), .ZN(n130) );
  INV_X1 U32 ( .A(n131), .ZN(Y[8]) );
  AOI22_X1 U33 ( .A1(A[8]), .A2(n67), .B1(B[8]), .B2(SEL), .ZN(n131) );
  INV_X1 U34 ( .A(n132), .ZN(Y[9]) );
  AOI22_X1 U35 ( .A1(A[9]), .A2(n67), .B1(SEL), .B2(B[9]), .ZN(n132) );
  INV_X1 U36 ( .A(n102), .ZN(Y[10]) );
  AOI22_X1 U37 ( .A1(A[10]), .A2(n33), .B1(B[10]), .B2(SEL), .ZN(n102) );
  INV_X1 U38 ( .A(n103), .ZN(Y[11]) );
  AOI22_X1 U39 ( .A1(A[11]), .A2(n33), .B1(B[11]), .B2(SEL), .ZN(n103) );
  INV_X1 U40 ( .A(n104), .ZN(Y[12]) );
  AOI22_X1 U41 ( .A1(A[12]), .A2(n33), .B1(B[12]), .B2(SEL), .ZN(n104) );
  INV_X1 U42 ( .A(n105), .ZN(Y[13]) );
  AOI22_X1 U43 ( .A1(A[13]), .A2(n33), .B1(B[13]), .B2(SEL), .ZN(n105) );
  INV_X1 U44 ( .A(n106), .ZN(Y[14]) );
  AOI22_X1 U45 ( .A1(A[14]), .A2(n33), .B1(B[14]), .B2(SEL), .ZN(n106) );
  INV_X1 U46 ( .A(n107), .ZN(Y[15]) );
  AOI22_X1 U47 ( .A1(A[15]), .A2(n33), .B1(B[15]), .B2(SEL), .ZN(n107) );
  INV_X1 U48 ( .A(n108), .ZN(Y[16]) );
  AOI22_X1 U49 ( .A1(A[16]), .A2(n33), .B1(B[16]), .B2(SEL), .ZN(n108) );
  INV_X1 U50 ( .A(n109), .ZN(Y[17]) );
  AOI22_X1 U51 ( .A1(A[17]), .A2(n33), .B1(B[17]), .B2(SEL), .ZN(n109) );
  INV_X1 U52 ( .A(n110), .ZN(Y[18]) );
  AOI22_X1 U53 ( .A1(A[18]), .A2(n33), .B1(B[18]), .B2(SEL), .ZN(n110) );
  INV_X1 U54 ( .A(n111), .ZN(Y[19]) );
  AOI22_X1 U55 ( .A1(A[19]), .A2(n33), .B1(B[19]), .B2(SEL), .ZN(n111) );
  INV_X1 U56 ( .A(n113), .ZN(Y[20]) );
  AOI22_X1 U57 ( .A1(A[20]), .A2(n66), .B1(B[20]), .B2(SEL), .ZN(n113) );
  INV_X1 U58 ( .A(n114), .ZN(Y[21]) );
  AOI22_X1 U59 ( .A1(A[21]), .A2(n66), .B1(B[21]), .B2(SEL), .ZN(n114) );
  INV_X1 U60 ( .A(n115), .ZN(Y[22]) );
  AOI22_X1 U61 ( .A1(A[22]), .A2(n66), .B1(B[22]), .B2(SEL), .ZN(n115) );
  INV_X1 U62 ( .A(n122), .ZN(Y[29]) );
  AOI22_X1 U63 ( .A1(A[29]), .A2(n66), .B1(B[29]), .B2(SEL), .ZN(n122) );
  INV_X1 U64 ( .A(n124), .ZN(Y[30]) );
  AOI22_X1 U65 ( .A1(A[30]), .A2(n66), .B1(B[30]), .B2(SEL), .ZN(n124) );
  INV_X1 U66 ( .A(n125), .ZN(Y[31]) );
  AOI22_X1 U67 ( .A1(A[31]), .A2(n67), .B1(B[31]), .B2(SEL), .ZN(n125) );
  INV_X1 U68 ( .A(SEL), .ZN(n100) );
endmodule


module REG_GEN_NBIT32_3 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n47), .Q(Q[31]), .QN(n145) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n47), .Q(Q[30]), .QN(n144) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n47), .Q(Q[29]), .QN(n143) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n47), .Q(Q[28]), .QN(n142) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n47), .Q(Q[27]), .QN(n141) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n47), .Q(Q[26]), .QN(n140) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n47), .Q(Q[25]), .QN(n139) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n47), .Q(Q[24]), .QN(n138) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n47), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n47), .Q(Q[22]), .QN(n136) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n47), .Q(Q[21]), .QN(n135) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n47), .Q(Q[20]), .QN(n134) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n48), .Q(Q[19]), .QN(n133) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n48), .Q(Q[18]), .QN(n132) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n48), .Q(Q[17]), .QN(n131) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n48), .Q(Q[16]), .QN(n130) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n48), .Q(Q[15]), .QN(n129) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n48), .Q(Q[14]), .QN(n128) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n48), .Q(Q[13]), .QN(n127) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n48), .Q(Q[12]), .QN(n126) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n48), .Q(Q[11]), .QN(n125) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n48), .Q(Q[10]), .QN(n124) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n48), .Q(Q[9]), .QN(n123) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n48), .Q(Q[8]), .QN(n122) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n49), .Q(Q[7]), .QN(n121) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n49), .Q(Q[6]), .QN(n120) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n49), .Q(Q[5]), .QN(n119) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n49), .Q(Q[4]), .QN(n118) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n49), .Q(Q[3]), .QN(n117) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n49), .Q(Q[2]), .QN(n116) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n49), .Q(Q[1]), .QN(n115) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n49), .Q(Q[0]), .QN(n114) );
  INV_X1 U2 ( .A(n46), .ZN(n37) );
  INV_X1 U3 ( .A(n46), .ZN(n36) );
  BUF_X1 U4 ( .A(n35), .Z(n46) );
  BUF_X1 U5 ( .A(n34), .Z(n41) );
  BUF_X1 U6 ( .A(n34), .Z(n42) );
  BUF_X1 U7 ( .A(n35), .Z(n44) );
  BUF_X1 U8 ( .A(n33), .Z(n38) );
  BUF_X1 U9 ( .A(n33), .Z(n39) );
  BUF_X1 U10 ( .A(n33), .Z(n40) );
  BUF_X1 U11 ( .A(n34), .Z(n43) );
  BUF_X1 U12 ( .A(n35), .Z(n45) );
  BUF_X1 U13 ( .A(RESET_n), .Z(n48) );
  BUF_X1 U14 ( .A(RESET_n), .Z(n47) );
  BUF_X1 U15 ( .A(RESET_n), .Z(n49) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n35) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n33) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n34) );
  OAI22_X1 U19 ( .A1(n114), .A2(n37), .B1(n39), .B2(n113), .ZN(n32) );
  INV_X1 U20 ( .A(D[0]), .ZN(n113) );
  OAI22_X1 U21 ( .A1(n115), .A2(n36), .B1(n39), .B2(n112), .ZN(n31) );
  INV_X1 U22 ( .A(D[1]), .ZN(n112) );
  OAI22_X1 U23 ( .A1(n137), .A2(n37), .B1(n38), .B2(n58), .ZN(n9) );
  INV_X1 U24 ( .A(D[23]), .ZN(n58) );
  OAI22_X1 U25 ( .A1(n138), .A2(n36), .B1(n38), .B2(n57), .ZN(n8) );
  INV_X1 U26 ( .A(D[24]), .ZN(n57) );
  OAI22_X1 U27 ( .A1(n139), .A2(n37), .B1(n38), .B2(n56), .ZN(n7) );
  INV_X1 U28 ( .A(D[25]), .ZN(n56) );
  OAI22_X1 U29 ( .A1(n140), .A2(n36), .B1(n38), .B2(n55), .ZN(n6) );
  INV_X1 U30 ( .A(D[26]), .ZN(n55) );
  OAI22_X1 U31 ( .A1(n141), .A2(n37), .B1(n39), .B2(n54), .ZN(n5) );
  INV_X1 U32 ( .A(D[27]), .ZN(n54) );
  OAI22_X1 U33 ( .A1(n142), .A2(n36), .B1(n39), .B2(n53), .ZN(n4) );
  INV_X1 U34 ( .A(D[28]), .ZN(n53) );
  OAI22_X1 U35 ( .A1(n116), .A2(n37), .B1(n40), .B2(n111), .ZN(n30) );
  INV_X1 U36 ( .A(D[2]), .ZN(n111) );
  OAI22_X1 U37 ( .A1(n117), .A2(n37), .B1(n40), .B2(n110), .ZN(n29) );
  INV_X1 U38 ( .A(D[3]), .ZN(n110) );
  OAI22_X1 U39 ( .A1(n118), .A2(n37), .B1(n40), .B2(n109), .ZN(n28) );
  INV_X1 U40 ( .A(D[4]), .ZN(n109) );
  OAI22_X1 U41 ( .A1(n119), .A2(n37), .B1(n41), .B2(n108), .ZN(n27) );
  INV_X1 U42 ( .A(D[5]), .ZN(n108) );
  OAI22_X1 U43 ( .A1(n120), .A2(n37), .B1(n41), .B2(n107), .ZN(n26) );
  INV_X1 U44 ( .A(D[6]), .ZN(n107) );
  OAI22_X1 U45 ( .A1(n121), .A2(n37), .B1(n41), .B2(n106), .ZN(n25) );
  INV_X1 U46 ( .A(D[7]), .ZN(n106) );
  OAI22_X1 U47 ( .A1(n122), .A2(n37), .B1(n41), .B2(n105), .ZN(n24) );
  INV_X1 U48 ( .A(D[8]), .ZN(n105) );
  OAI22_X1 U49 ( .A1(n123), .A2(n37), .B1(n42), .B2(n104), .ZN(n23) );
  INV_X1 U50 ( .A(D[9]), .ZN(n104) );
  OAI22_X1 U51 ( .A1(n124), .A2(n37), .B1(n42), .B2(n103), .ZN(n22) );
  INV_X1 U52 ( .A(D[10]), .ZN(n103) );
  OAI22_X1 U53 ( .A1(n125), .A2(n37), .B1(n42), .B2(n102), .ZN(n21) );
  INV_X1 U54 ( .A(D[11]), .ZN(n102) );
  OAI22_X1 U55 ( .A1(n126), .A2(n37), .B1(n42), .B2(n101), .ZN(n20) );
  INV_X1 U56 ( .A(D[12]), .ZN(n101) );
  OAI22_X1 U57 ( .A1(n127), .A2(n36), .B1(n43), .B2(n100), .ZN(n19) );
  INV_X1 U58 ( .A(D[13]), .ZN(n100) );
  OAI22_X1 U59 ( .A1(n128), .A2(n36), .B1(n43), .B2(n99), .ZN(n18) );
  INV_X1 U60 ( .A(D[14]), .ZN(n99) );
  OAI22_X1 U61 ( .A1(n129), .A2(n36), .B1(n43), .B2(n98), .ZN(n17) );
  INV_X1 U62 ( .A(D[15]), .ZN(n98) );
  OAI22_X1 U63 ( .A1(n130), .A2(n36), .B1(n44), .B2(n65), .ZN(n16) );
  INV_X1 U64 ( .A(D[16]), .ZN(n65) );
  OAI22_X1 U65 ( .A1(n131), .A2(n36), .B1(n44), .B2(n64), .ZN(n15) );
  INV_X1 U66 ( .A(D[17]), .ZN(n64) );
  OAI22_X1 U67 ( .A1(n132), .A2(n36), .B1(n44), .B2(n63), .ZN(n14) );
  INV_X1 U68 ( .A(D[18]), .ZN(n63) );
  OAI22_X1 U69 ( .A1(n133), .A2(n36), .B1(n44), .B2(n62), .ZN(n13) );
  INV_X1 U70 ( .A(D[19]), .ZN(n62) );
  OAI22_X1 U71 ( .A1(n134), .A2(n36), .B1(n45), .B2(n61), .ZN(n12) );
  INV_X1 U72 ( .A(D[20]), .ZN(n61) );
  OAI22_X1 U73 ( .A1(n135), .A2(n36), .B1(n45), .B2(n60), .ZN(n11) );
  INV_X1 U74 ( .A(D[21]), .ZN(n60) );
  OAI22_X1 U75 ( .A1(n136), .A2(n36), .B1(n45), .B2(n59), .ZN(n10) );
  INV_X1 U76 ( .A(D[22]), .ZN(n59) );
  OAI22_X1 U77 ( .A1(n143), .A2(n37), .B1(n40), .B2(n52), .ZN(n3) );
  INV_X1 U78 ( .A(D[29]), .ZN(n52) );
  OAI22_X1 U79 ( .A1(n144), .A2(n36), .B1(n43), .B2(n51), .ZN(n2) );
  INV_X1 U80 ( .A(D[30]), .ZN(n51) );
  OAI22_X1 U81 ( .A1(n145), .A2(n36), .B1(n45), .B2(n50), .ZN(n1) );
  INV_X1 U82 ( .A(D[31]), .ZN(n50) );
endmodule


module REG_GEN_NBIT32_2 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n49), .Q(Q[31]), .QN(n145) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n49), .Q(Q[30]), .QN(n144) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n49), .Q(Q[29]), .QN(n143) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n49), .Q(Q[28]), .QN(n142) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n49), .Q(Q[27]), .QN(n141) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n49), .Q(Q[26]), .QN(n140) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n49), .Q(Q[25]), .QN(n139) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n49), .Q(Q[24]), .QN(n138) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n48), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n48), .Q(Q[22]), .QN(n136) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n48), .Q(Q[21]), .QN(n135) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n48), .Q(Q[20]), .QN(n134) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n48), .Q(Q[19]), .QN(n133) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n48), .Q(Q[18]), .QN(n132) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n48), .Q(Q[17]), .QN(n131) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n48), .Q(Q[16]), .QN(n130) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n48), .Q(Q[15]), .QN(n129) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n48), .Q(Q[14]), .QN(n128) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n48), .Q(Q[13]), .QN(n127) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n48), .Q(Q[12]), .QN(n126) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n47), .Q(Q[11]), .QN(n125) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n47), .Q(Q[10]), .QN(n124) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n47), .Q(Q[9]), .QN(n123) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n47), .Q(Q[8]), .QN(n122) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n47), .Q(Q[7]), .QN(n121) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n47), .Q(Q[6]), .QN(n120) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n47), .Q(Q[5]), .QN(n119) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n47), .Q(Q[4]), .QN(n118) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n47), .Q(Q[3]), .QN(n117) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n47), .Q(Q[2]), .QN(n116) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n47), .Q(Q[1]), .QN(n115) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n47), .Q(Q[0]), .QN(n114) );
  INV_X1 U2 ( .A(n46), .ZN(n37) );
  INV_X1 U3 ( .A(n46), .ZN(n36) );
  BUF_X1 U4 ( .A(n35), .Z(n46) );
  BUF_X1 U5 ( .A(n34), .Z(n41) );
  BUF_X1 U6 ( .A(n34), .Z(n42) );
  BUF_X1 U7 ( .A(n35), .Z(n44) );
  BUF_X1 U8 ( .A(n33), .Z(n38) );
  BUF_X1 U9 ( .A(n33), .Z(n39) );
  BUF_X1 U10 ( .A(n33), .Z(n40) );
  BUF_X1 U11 ( .A(n34), .Z(n43) );
  BUF_X1 U12 ( .A(n35), .Z(n45) );
  BUF_X1 U13 ( .A(RESET_n), .Z(n47) );
  BUF_X1 U14 ( .A(RESET_n), .Z(n48) );
  BUF_X1 U15 ( .A(RESET_n), .Z(n49) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n35) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n33) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n34) );
  OAI22_X1 U19 ( .A1(n114), .A2(n37), .B1(n39), .B2(n113), .ZN(n32) );
  INV_X1 U20 ( .A(D[0]), .ZN(n113) );
  OAI22_X1 U21 ( .A1(n115), .A2(n36), .B1(n39), .B2(n112), .ZN(n31) );
  INV_X1 U22 ( .A(D[1]), .ZN(n112) );
  OAI22_X1 U23 ( .A1(n137), .A2(n37), .B1(n38), .B2(n58), .ZN(n9) );
  INV_X1 U24 ( .A(D[23]), .ZN(n58) );
  OAI22_X1 U25 ( .A1(n138), .A2(n36), .B1(n38), .B2(n57), .ZN(n8) );
  INV_X1 U26 ( .A(D[24]), .ZN(n57) );
  OAI22_X1 U27 ( .A1(n139), .A2(n37), .B1(n38), .B2(n56), .ZN(n7) );
  INV_X1 U28 ( .A(D[25]), .ZN(n56) );
  OAI22_X1 U29 ( .A1(n140), .A2(n36), .B1(n38), .B2(n55), .ZN(n6) );
  INV_X1 U30 ( .A(D[26]), .ZN(n55) );
  OAI22_X1 U31 ( .A1(n141), .A2(n37), .B1(n39), .B2(n54), .ZN(n5) );
  INV_X1 U32 ( .A(D[27]), .ZN(n54) );
  OAI22_X1 U33 ( .A1(n142), .A2(n36), .B1(n39), .B2(n53), .ZN(n4) );
  INV_X1 U34 ( .A(D[28]), .ZN(n53) );
  OAI22_X1 U35 ( .A1(n116), .A2(n37), .B1(n40), .B2(n111), .ZN(n30) );
  INV_X1 U36 ( .A(D[2]), .ZN(n111) );
  OAI22_X1 U37 ( .A1(n117), .A2(n37), .B1(n40), .B2(n110), .ZN(n29) );
  INV_X1 U38 ( .A(D[3]), .ZN(n110) );
  OAI22_X1 U39 ( .A1(n118), .A2(n37), .B1(n40), .B2(n109), .ZN(n28) );
  INV_X1 U40 ( .A(D[4]), .ZN(n109) );
  OAI22_X1 U41 ( .A1(n119), .A2(n37), .B1(n41), .B2(n108), .ZN(n27) );
  INV_X1 U42 ( .A(D[5]), .ZN(n108) );
  OAI22_X1 U43 ( .A1(n120), .A2(n37), .B1(n41), .B2(n107), .ZN(n26) );
  INV_X1 U44 ( .A(D[6]), .ZN(n107) );
  OAI22_X1 U45 ( .A1(n121), .A2(n37), .B1(n41), .B2(n106), .ZN(n25) );
  INV_X1 U46 ( .A(D[7]), .ZN(n106) );
  OAI22_X1 U47 ( .A1(n122), .A2(n37), .B1(n41), .B2(n105), .ZN(n24) );
  INV_X1 U48 ( .A(D[8]), .ZN(n105) );
  OAI22_X1 U49 ( .A1(n123), .A2(n37), .B1(n42), .B2(n104), .ZN(n23) );
  INV_X1 U50 ( .A(D[9]), .ZN(n104) );
  OAI22_X1 U51 ( .A1(n124), .A2(n37), .B1(n42), .B2(n103), .ZN(n22) );
  INV_X1 U52 ( .A(D[10]), .ZN(n103) );
  OAI22_X1 U53 ( .A1(n125), .A2(n37), .B1(n42), .B2(n102), .ZN(n21) );
  INV_X1 U54 ( .A(D[11]), .ZN(n102) );
  OAI22_X1 U55 ( .A1(n126), .A2(n37), .B1(n42), .B2(n101), .ZN(n20) );
  INV_X1 U56 ( .A(D[12]), .ZN(n101) );
  OAI22_X1 U57 ( .A1(n127), .A2(n36), .B1(n43), .B2(n100), .ZN(n19) );
  INV_X1 U58 ( .A(D[13]), .ZN(n100) );
  OAI22_X1 U59 ( .A1(n128), .A2(n36), .B1(n43), .B2(n99), .ZN(n18) );
  INV_X1 U60 ( .A(D[14]), .ZN(n99) );
  OAI22_X1 U61 ( .A1(n129), .A2(n36), .B1(n43), .B2(n98), .ZN(n17) );
  INV_X1 U62 ( .A(D[15]), .ZN(n98) );
  OAI22_X1 U63 ( .A1(n130), .A2(n36), .B1(n44), .B2(n65), .ZN(n16) );
  INV_X1 U64 ( .A(D[16]), .ZN(n65) );
  OAI22_X1 U65 ( .A1(n131), .A2(n36), .B1(n44), .B2(n64), .ZN(n15) );
  INV_X1 U66 ( .A(D[17]), .ZN(n64) );
  OAI22_X1 U67 ( .A1(n132), .A2(n36), .B1(n44), .B2(n63), .ZN(n14) );
  INV_X1 U68 ( .A(D[18]), .ZN(n63) );
  OAI22_X1 U69 ( .A1(n133), .A2(n36), .B1(n44), .B2(n62), .ZN(n13) );
  INV_X1 U70 ( .A(D[19]), .ZN(n62) );
  OAI22_X1 U71 ( .A1(n134), .A2(n36), .B1(n45), .B2(n61), .ZN(n12) );
  INV_X1 U72 ( .A(D[20]), .ZN(n61) );
  OAI22_X1 U73 ( .A1(n135), .A2(n36), .B1(n45), .B2(n60), .ZN(n11) );
  INV_X1 U74 ( .A(D[21]), .ZN(n60) );
  OAI22_X1 U75 ( .A1(n136), .A2(n36), .B1(n45), .B2(n59), .ZN(n10) );
  INV_X1 U76 ( .A(D[22]), .ZN(n59) );
  OAI22_X1 U77 ( .A1(n143), .A2(n37), .B1(n40), .B2(n52), .ZN(n3) );
  INV_X1 U78 ( .A(D[29]), .ZN(n52) );
  OAI22_X1 U79 ( .A1(n144), .A2(n36), .B1(n43), .B2(n51), .ZN(n2) );
  INV_X1 U80 ( .A(D[30]), .ZN(n51) );
  OAI22_X1 U81 ( .A1(n145), .A2(n36), .B1(n45), .B2(n50), .ZN(n1) );
  INV_X1 U82 ( .A(D[31]), .ZN(n50) );
endmodule


module REG_GEN_NBIT32_1 ( D, CK, Enable_n, RESET_n, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, Enable_n, RESET_n;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n47), .Q(Q[31]), .QN(n66) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n49), .Q(Q[30]), .QN(n67) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n49), .Q(Q[29]), .QN(n68) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n49), .Q(Q[28]), .QN(n69) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n49), .Q(Q[27]), .QN(n70) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n48), .Q(Q[26]), .QN(n71) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n49), .Q(Q[25]), .QN(n72) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n48), .Q(Q[24]), .QN(n73) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n48), .Q(Q[23]), .QN(n74) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n48), .Q(Q[22]), .QN(n75) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n48), .Q(Q[21]), .QN(n76) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n49), .Q(Q[20]), .QN(n77) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n48), .Q(Q[19]), .QN(n78) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n48), .Q(Q[18]), .QN(n79) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n49), .Q(Q[17]), .QN(n80) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n48), .Q(Q[16]), .QN(n81) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n48), .Q(Q[15]), .QN(n82) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n48), .Q(Q[14]), .QN(n83) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n47), .Q(Q[13]), .QN(n84) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n48), .Q(Q[12]), .QN(n85) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n47), .Q(Q[11]), .QN(n86) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n47), .Q(Q[10]), .QN(n87) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n47), .Q(Q[9]), .QN(n88) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n47), .Q(Q[8]), .QN(n89) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n47), .Q(Q[7]), .QN(n90) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n47), .Q(Q[6]), .QN(n91) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n47), .Q(Q[5]), .QN(n92) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n47), .Q(Q[4]), .QN(n93) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n47), .Q(Q[3]), .QN(n94) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n47), .Q(Q[2]), .QN(n95) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n48), .Q(Q[1]), .QN(n96) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n49), .Q(Q[0]), .QN(n97) );
  INV_X1 U2 ( .A(n46), .ZN(n37) );
  INV_X1 U3 ( .A(n46), .ZN(n36) );
  BUF_X1 U4 ( .A(n35), .Z(n46) );
  BUF_X1 U5 ( .A(n34), .Z(n41) );
  BUF_X1 U6 ( .A(n34), .Z(n42) );
  BUF_X1 U7 ( .A(n35), .Z(n44) );
  BUF_X1 U8 ( .A(n33), .Z(n38) );
  BUF_X1 U9 ( .A(n33), .Z(n39) );
  BUF_X1 U10 ( .A(n33), .Z(n40) );
  BUF_X1 U11 ( .A(n34), .Z(n43) );
  BUF_X1 U12 ( .A(n35), .Z(n45) );
  BUF_X1 U13 ( .A(RESET_n), .Z(n48) );
  BUF_X1 U14 ( .A(RESET_n), .Z(n47) );
  BUF_X1 U15 ( .A(RESET_n), .Z(n49) );
  BUF_X1 U16 ( .A(Enable_n), .Z(n35) );
  BUF_X1 U17 ( .A(Enable_n), .Z(n33) );
  BUF_X1 U18 ( .A(Enable_n), .Z(n34) );
  OAI22_X1 U19 ( .A1(n70), .A2(n37), .B1(n39), .B2(n54), .ZN(n5) );
  INV_X1 U20 ( .A(D[27]), .ZN(n54) );
  OAI22_X1 U21 ( .A1(n69), .A2(n36), .B1(n39), .B2(n53), .ZN(n4) );
  INV_X1 U22 ( .A(D[28]), .ZN(n53) );
  OAI22_X1 U23 ( .A1(n97), .A2(n37), .B1(n39), .B2(n113), .ZN(n32) );
  INV_X1 U24 ( .A(D[0]), .ZN(n113) );
  OAI22_X1 U25 ( .A1(n96), .A2(n36), .B1(n39), .B2(n112), .ZN(n31) );
  INV_X1 U26 ( .A(D[1]), .ZN(n112) );
  OAI22_X1 U27 ( .A1(n74), .A2(n37), .B1(n38), .B2(n58), .ZN(n9) );
  INV_X1 U28 ( .A(D[23]), .ZN(n58) );
  OAI22_X1 U29 ( .A1(n73), .A2(n36), .B1(n38), .B2(n57), .ZN(n8) );
  INV_X1 U30 ( .A(D[24]), .ZN(n57) );
  OAI22_X1 U31 ( .A1(n72), .A2(n37), .B1(n38), .B2(n56), .ZN(n7) );
  INV_X1 U32 ( .A(D[25]), .ZN(n56) );
  OAI22_X1 U33 ( .A1(n71), .A2(n36), .B1(n38), .B2(n55), .ZN(n6) );
  INV_X1 U34 ( .A(D[26]), .ZN(n55) );
  OAI22_X1 U35 ( .A1(n95), .A2(n37), .B1(n40), .B2(n111), .ZN(n30) );
  INV_X1 U36 ( .A(D[2]), .ZN(n111) );
  OAI22_X1 U37 ( .A1(n94), .A2(n37), .B1(n40), .B2(n110), .ZN(n29) );
  INV_X1 U38 ( .A(D[3]), .ZN(n110) );
  OAI22_X1 U39 ( .A1(n93), .A2(n37), .B1(n40), .B2(n109), .ZN(n28) );
  INV_X1 U40 ( .A(D[4]), .ZN(n109) );
  OAI22_X1 U41 ( .A1(n92), .A2(n37), .B1(n41), .B2(n108), .ZN(n27) );
  INV_X1 U42 ( .A(D[5]), .ZN(n108) );
  OAI22_X1 U43 ( .A1(n91), .A2(n37), .B1(n41), .B2(n107), .ZN(n26) );
  INV_X1 U44 ( .A(D[6]), .ZN(n107) );
  OAI22_X1 U45 ( .A1(n90), .A2(n37), .B1(n41), .B2(n106), .ZN(n25) );
  INV_X1 U46 ( .A(D[7]), .ZN(n106) );
  OAI22_X1 U47 ( .A1(n89), .A2(n37), .B1(n41), .B2(n105), .ZN(n24) );
  INV_X1 U48 ( .A(D[8]), .ZN(n105) );
  OAI22_X1 U49 ( .A1(n88), .A2(n37), .B1(n42), .B2(n104), .ZN(n23) );
  INV_X1 U50 ( .A(D[9]), .ZN(n104) );
  OAI22_X1 U51 ( .A1(n87), .A2(n37), .B1(n42), .B2(n103), .ZN(n22) );
  INV_X1 U52 ( .A(D[10]), .ZN(n103) );
  OAI22_X1 U53 ( .A1(n86), .A2(n37), .B1(n42), .B2(n102), .ZN(n21) );
  INV_X1 U54 ( .A(D[11]), .ZN(n102) );
  OAI22_X1 U55 ( .A1(n85), .A2(n37), .B1(n42), .B2(n101), .ZN(n20) );
  INV_X1 U56 ( .A(D[12]), .ZN(n101) );
  OAI22_X1 U57 ( .A1(n84), .A2(n36), .B1(n43), .B2(n100), .ZN(n19) );
  INV_X1 U58 ( .A(D[13]), .ZN(n100) );
  OAI22_X1 U59 ( .A1(n83), .A2(n36), .B1(n43), .B2(n99), .ZN(n18) );
  INV_X1 U60 ( .A(D[14]), .ZN(n99) );
  OAI22_X1 U61 ( .A1(n82), .A2(n36), .B1(n43), .B2(n98), .ZN(n17) );
  INV_X1 U62 ( .A(D[15]), .ZN(n98) );
  OAI22_X1 U63 ( .A1(n81), .A2(n36), .B1(n44), .B2(n65), .ZN(n16) );
  INV_X1 U64 ( .A(D[16]), .ZN(n65) );
  OAI22_X1 U65 ( .A1(n80), .A2(n36), .B1(n44), .B2(n64), .ZN(n15) );
  INV_X1 U66 ( .A(D[17]), .ZN(n64) );
  OAI22_X1 U67 ( .A1(n79), .A2(n36), .B1(n44), .B2(n63), .ZN(n14) );
  INV_X1 U68 ( .A(D[18]), .ZN(n63) );
  OAI22_X1 U69 ( .A1(n78), .A2(n36), .B1(n44), .B2(n62), .ZN(n13) );
  INV_X1 U70 ( .A(D[19]), .ZN(n62) );
  OAI22_X1 U71 ( .A1(n77), .A2(n36), .B1(n45), .B2(n61), .ZN(n12) );
  INV_X1 U72 ( .A(D[20]), .ZN(n61) );
  OAI22_X1 U73 ( .A1(n76), .A2(n36), .B1(n45), .B2(n60), .ZN(n11) );
  INV_X1 U74 ( .A(D[21]), .ZN(n60) );
  OAI22_X1 U75 ( .A1(n75), .A2(n36), .B1(n45), .B2(n59), .ZN(n10) );
  INV_X1 U76 ( .A(D[22]), .ZN(n59) );
  OAI22_X1 U77 ( .A1(n68), .A2(n37), .B1(n40), .B2(n52), .ZN(n3) );
  INV_X1 U78 ( .A(D[29]), .ZN(n52) );
  OAI22_X1 U79 ( .A1(n67), .A2(n36), .B1(n43), .B2(n51), .ZN(n2) );
  INV_X1 U80 ( .A(D[30]), .ZN(n51) );
  OAI22_X1 U81 ( .A1(n66), .A2(n36), .B1(n45), .B2(n50), .ZN(n1) );
  INV_X1 U82 ( .A(D[31]), .ZN(n50) );
endmodule


module memoryUnit_nbit32 ( rst, clk, en_reg, b_op, j_op, jal_op, alu_out, 
        r2_out, PC, lab_b, lab_j, rw_exe, dataout_from_mem, addr_mem, 
        datain_mem, next_PC, alu_out_mem, rw_mem, data_out );
  input [31:0] alu_out;
  input [31:0] r2_out;
  input [31:0] PC;
  input [31:0] lab_b;
  input [31:0] lab_j;
  input [31:0] rw_exe;
  input [31:0] dataout_from_mem;
  output [31:0] addr_mem;
  output [31:0] datain_mem;
  output [31:0] next_PC;
  output [31:0] alu_out_mem;
  output [31:0] rw_mem;
  output [31:0] data_out;
  input rst, clk, en_reg, b_op, j_op, jal_op;

  wire   [31:0] branch_pc;
  wire   [31:0] rf_out;
  wire   [31:0] rw_out;
  assign addr_mem[31] = alu_out[31];
  assign addr_mem[30] = alu_out[30];
  assign addr_mem[29] = alu_out[29];
  assign addr_mem[28] = alu_out[28];
  assign addr_mem[27] = alu_out[27];
  assign addr_mem[26] = alu_out[26];
  assign addr_mem[25] = alu_out[25];
  assign addr_mem[24] = alu_out[24];
  assign addr_mem[23] = alu_out[23];
  assign addr_mem[22] = alu_out[22];
  assign addr_mem[21] = alu_out[21];
  assign addr_mem[20] = alu_out[20];
  assign addr_mem[19] = alu_out[19];
  assign addr_mem[18] = alu_out[18];
  assign addr_mem[17] = alu_out[17];
  assign addr_mem[16] = alu_out[16];
  assign addr_mem[15] = alu_out[15];
  assign addr_mem[14] = alu_out[14];
  assign addr_mem[13] = alu_out[13];
  assign addr_mem[12] = alu_out[12];
  assign addr_mem[11] = alu_out[11];
  assign addr_mem[10] = alu_out[10];
  assign addr_mem[9] = alu_out[9];
  assign addr_mem[8] = alu_out[8];
  assign addr_mem[7] = alu_out[7];
  assign addr_mem[6] = alu_out[6];
  assign addr_mem[5] = alu_out[5];
  assign addr_mem[4] = alu_out[4];
  assign addr_mem[3] = alu_out[3];
  assign addr_mem[2] = alu_out[2];
  assign addr_mem[1] = alu_out[1];
  assign addr_mem[0] = alu_out[0];
  assign datain_mem[31] = r2_out[31];
  assign datain_mem[30] = r2_out[30];
  assign datain_mem[29] = r2_out[29];
  assign datain_mem[28] = r2_out[28];
  assign datain_mem[27] = r2_out[27];
  assign datain_mem[26] = r2_out[26];
  assign datain_mem[25] = r2_out[25];
  assign datain_mem[24] = r2_out[24];
  assign datain_mem[23] = r2_out[23];
  assign datain_mem[22] = r2_out[22];
  assign datain_mem[21] = r2_out[21];
  assign datain_mem[20] = r2_out[20];
  assign datain_mem[19] = r2_out[19];
  assign datain_mem[18] = r2_out[18];
  assign datain_mem[17] = r2_out[17];
  assign datain_mem[16] = r2_out[16];
  assign datain_mem[15] = r2_out[15];
  assign datain_mem[14] = r2_out[14];
  assign datain_mem[13] = r2_out[13];
  assign datain_mem[12] = r2_out[12];
  assign datain_mem[11] = r2_out[11];
  assign datain_mem[10] = r2_out[10];
  assign datain_mem[9] = r2_out[9];
  assign datain_mem[8] = r2_out[8];
  assign datain_mem[7] = r2_out[7];
  assign datain_mem[6] = r2_out[6];
  assign datain_mem[5] = r2_out[5];
  assign datain_mem[4] = r2_out[4];
  assign datain_mem[3] = r2_out[3];
  assign datain_mem[2] = r2_out[2];
  assign datain_mem[1] = r2_out[1];
  assign datain_mem[0] = r2_out[0];

  branch_block_nbit32 br_unit ( .branch_op(b_op), .cmp_out(alu_out), .PC(PC), 
        .label_PC(lab_b), .next_PC(branch_pc) );
  MUX21_GENERIC_NBIT32_6 jmp_unit ( .A(branch_pc), .B(lab_j), .SEL(j_op), .Y(
        next_PC) );
  MUX21_GENERIC_NBIT32_5 mux_jal_pc ( .A(dataout_from_mem), .B(PC), .SEL(
        jal_op), .Y(rf_out) );
  MUX21_GENERIC_NBIT32_4 mux_jal_r31 ( .A(rw_exe), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(jal_op), .Y(rw_out) );
  REG_GEN_NBIT32_3 mem_reg ( .D(rf_out), .CK(clk), .Enable_n(en_reg), 
        .RESET_n(rst), .Q(data_out) );
  REG_GEN_NBIT32_2 rw_reg ( .D(rw_out), .CK(clk), .Enable_n(en_reg), .RESET_n(
        rst), .Q(rw_mem) );
  REG_GEN_NBIT32_1 alu_reg ( .D(alu_out), .CK(clk), .Enable_n(en_reg), 
        .RESET_n(rst), .Q(alu_out_mem) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n33, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142;

  INV_X1 U1 ( .A(n78), .ZN(n68) );
  INV_X1 U2 ( .A(n78), .ZN(n69) );
  BUF_X1 U3 ( .A(n33), .Z(n70) );
  BUF_X1 U4 ( .A(n67), .Z(n76) );
  BUF_X1 U5 ( .A(n66), .Z(n75) );
  BUF_X1 U6 ( .A(n66), .Z(n73) );
  BUF_X1 U7 ( .A(n33), .Z(n72) );
  BUF_X1 U8 ( .A(n66), .Z(n74) );
  BUF_X1 U9 ( .A(n33), .Z(n71) );
  BUF_X1 U10 ( .A(n67), .Z(n78) );
  BUF_X1 U11 ( .A(n67), .Z(n77) );
  BUF_X1 U12 ( .A(SEL), .Z(n67) );
  BUF_X1 U13 ( .A(SEL), .Z(n66) );
  BUF_X1 U14 ( .A(SEL), .Z(n33) );
  INV_X1 U15 ( .A(n136), .ZN(Y[3]) );
  AOI22_X1 U16 ( .A1(A[3]), .A2(n68), .B1(B[3]), .B2(n71), .ZN(n136) );
  INV_X1 U17 ( .A(n137), .ZN(Y[4]) );
  AOI22_X1 U18 ( .A1(A[4]), .A2(n69), .B1(B[4]), .B2(n71), .ZN(n137) );
  INV_X1 U19 ( .A(n138), .ZN(Y[5]) );
  AOI22_X1 U20 ( .A1(A[5]), .A2(n68), .B1(B[5]), .B2(n70), .ZN(n138) );
  INV_X1 U21 ( .A(n139), .ZN(Y[6]) );
  AOI22_X1 U22 ( .A1(A[6]), .A2(n69), .B1(B[6]), .B2(n70), .ZN(n139) );
  INV_X1 U23 ( .A(n140), .ZN(Y[7]) );
  AOI22_X1 U24 ( .A1(A[7]), .A2(n68), .B1(B[7]), .B2(n70), .ZN(n140) );
  INV_X1 U25 ( .A(n141), .ZN(Y[8]) );
  AOI22_X1 U26 ( .A1(A[8]), .A2(n69), .B1(B[8]), .B2(n70), .ZN(n141) );
  INV_X1 U27 ( .A(n142), .ZN(Y[9]) );
  AOI22_X1 U28 ( .A1(A[9]), .A2(n68), .B1(n77), .B2(B[9]), .ZN(n142) );
  INV_X1 U29 ( .A(n135), .ZN(Y[31]) );
  AOI22_X1 U30 ( .A1(A[31]), .A2(n69), .B1(B[31]), .B2(n71), .ZN(n135) );
  INV_X1 U31 ( .A(n111), .ZN(Y[0]) );
  AOI22_X1 U32 ( .A1(A[0]), .A2(n68), .B1(B[0]), .B2(n77), .ZN(n111) );
  INV_X1 U33 ( .A(n122), .ZN(Y[1]) );
  AOI22_X1 U34 ( .A1(A[1]), .A2(n68), .B1(B[1]), .B2(n74), .ZN(n122) );
  INV_X1 U35 ( .A(n133), .ZN(Y[2]) );
  AOI22_X1 U36 ( .A1(A[2]), .A2(n69), .B1(B[2]), .B2(n71), .ZN(n133) );
  INV_X1 U37 ( .A(n112), .ZN(Y[10]) );
  AOI22_X1 U38 ( .A1(A[10]), .A2(n68), .B1(B[10]), .B2(n77), .ZN(n112) );
  INV_X1 U39 ( .A(n113), .ZN(Y[11]) );
  AOI22_X1 U40 ( .A1(A[11]), .A2(n68), .B1(B[11]), .B2(n77), .ZN(n113) );
  INV_X1 U41 ( .A(n114), .ZN(Y[12]) );
  AOI22_X1 U42 ( .A1(A[12]), .A2(n68), .B1(B[12]), .B2(n76), .ZN(n114) );
  INV_X1 U43 ( .A(n115), .ZN(Y[13]) );
  AOI22_X1 U44 ( .A1(A[13]), .A2(n68), .B1(B[13]), .B2(n76), .ZN(n115) );
  INV_X1 U45 ( .A(n116), .ZN(Y[14]) );
  AOI22_X1 U46 ( .A1(A[14]), .A2(n68), .B1(B[14]), .B2(n76), .ZN(n116) );
  INV_X1 U47 ( .A(n117), .ZN(Y[15]) );
  AOI22_X1 U48 ( .A1(A[15]), .A2(n68), .B1(B[15]), .B2(n76), .ZN(n117) );
  INV_X1 U49 ( .A(n118), .ZN(Y[16]) );
  AOI22_X1 U50 ( .A1(A[16]), .A2(n68), .B1(B[16]), .B2(n75), .ZN(n118) );
  INV_X1 U51 ( .A(n119), .ZN(Y[17]) );
  AOI22_X1 U52 ( .A1(A[17]), .A2(n68), .B1(B[17]), .B2(n75), .ZN(n119) );
  INV_X1 U53 ( .A(n120), .ZN(Y[18]) );
  AOI22_X1 U54 ( .A1(A[18]), .A2(n68), .B1(B[18]), .B2(n75), .ZN(n120) );
  INV_X1 U55 ( .A(n121), .ZN(Y[19]) );
  AOI22_X1 U56 ( .A1(A[19]), .A2(n68), .B1(B[19]), .B2(n75), .ZN(n121) );
  INV_X1 U57 ( .A(n123), .ZN(Y[20]) );
  AOI22_X1 U58 ( .A1(A[20]), .A2(n69), .B1(B[20]), .B2(n74), .ZN(n123) );
  INV_X1 U59 ( .A(n124), .ZN(Y[21]) );
  AOI22_X1 U60 ( .A1(A[21]), .A2(n69), .B1(B[21]), .B2(n74), .ZN(n124) );
  INV_X1 U61 ( .A(n125), .ZN(Y[22]) );
  AOI22_X1 U62 ( .A1(A[22]), .A2(n69), .B1(B[22]), .B2(n73), .ZN(n125) );
  INV_X1 U63 ( .A(n126), .ZN(Y[23]) );
  AOI22_X1 U64 ( .A1(A[23]), .A2(n69), .B1(B[23]), .B2(n73), .ZN(n126) );
  INV_X1 U65 ( .A(n127), .ZN(Y[24]) );
  AOI22_X1 U66 ( .A1(A[24]), .A2(n69), .B1(B[24]), .B2(n73), .ZN(n127) );
  INV_X1 U67 ( .A(n128), .ZN(Y[25]) );
  AOI22_X1 U68 ( .A1(A[25]), .A2(n69), .B1(B[25]), .B2(n73), .ZN(n128) );
  INV_X1 U69 ( .A(n129), .ZN(Y[26]) );
  AOI22_X1 U70 ( .A1(A[26]), .A2(n69), .B1(B[26]), .B2(n72), .ZN(n129) );
  INV_X1 U71 ( .A(n130), .ZN(Y[27]) );
  AOI22_X1 U72 ( .A1(A[27]), .A2(n69), .B1(B[27]), .B2(n72), .ZN(n130) );
  INV_X1 U73 ( .A(n131), .ZN(Y[28]) );
  AOI22_X1 U74 ( .A1(A[28]), .A2(n69), .B1(B[28]), .B2(n72), .ZN(n131) );
  INV_X1 U75 ( .A(n132), .ZN(Y[29]) );
  AOI22_X1 U76 ( .A1(A[29]), .A2(n69), .B1(B[29]), .B2(n72), .ZN(n132) );
  INV_X1 U77 ( .A(n134), .ZN(Y[30]) );
  AOI22_X1 U78 ( .A1(A[30]), .A2(n69), .B1(B[30]), .B2(n74), .ZN(n134) );
endmodule


module writeBackUnit_nbit32 ( MemtoReg, ReadData, AluResult, WriteData );
  input [31:0] ReadData;
  input [31:0] AluResult;
  output [31:0] WriteData;
  input MemtoReg;


  MUX21_GENERIC_NBIT32_3 mux_writeBack ( .A(ReadData), .B(AluResult), .SEL(
        MemtoReg), .Y(WriteData) );
endmodule


module datapath_nbit32 ( Clk, Rst, PC_op, en_reg_if, RD1, RD2, dout_IRAM, 
        addr_IRAM, en_reg_id, WR, Opcode, Func, sel_ex, sel_mux_rw, en_reg_ex, 
        alu_sel, en_reg_mem, dataout_from_mem, addr_mem, datain_mem, b_op_mem, 
        j_op_mem, jal_op_mem, MemtoReg_wb, pipe_out );
  input [31:0] dout_IRAM;
  output [31:0] addr_IRAM;
  output [5:0] Opcode;
  output [10:0] Func;
  input [3:0] alu_sel;
  input [31:0] dataout_from_mem;
  output [31:0] addr_mem;
  output [31:0] datain_mem;
  output [31:0] pipe_out;
  input Clk, Rst, PC_op, en_reg_if, RD1, RD2, en_reg_id, WR, sel_ex,
         sel_mux_rw, en_reg_ex, en_reg_mem, b_op_mem, j_op_mem, jal_op_mem,
         MemtoReg_wb;
  wire   n1;
  wire   [31:0] pc_from_mem_to_fetch;
  wire   [31:0] PC_Next_fetch;
  wire   [31:0] IRAM;
  wire   [4:0] ADD_RW;
  wire   [31:0] RW_R_decode;
  wire   [31:0] RW_I_decode;
  wire   [31:0] J_imm;
  wire   [31:0] I_imm;
  wire   [31:0] RD_data_1;
  wire   [31:0] RD_data_2;
  wire   [31:0] PC_Next_decode;
  wire   [31:0] alu_out;
  wire   [31:0] aluR2_to_mem;
  wire   [31:0] b_from_ex_to_mem;
  wire   [31:0] pc_from_ex_to_mem;
  wire   [31:0] rw_from_ex_to_mem;
  wire   [31:0] j_from_ex_to_mem;
  wire   [31:0] alu_out_mem;
  wire   [31:0] data_from_mem_to_wb;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26;

  fetchUnit_nbit32 IFU ( .Clk(Clk), .Rst(n1), .en_reg(en_reg_if), 
        .PC_branch_jump(pc_from_mem_to_fetch), .dout_IRAM(dout_IRAM), .PC_op(
        PC_op), .PC_Next_out(PC_Next_fetch), .addr_IRAM(addr_IRAM), 
        .IRAM_reg_out(IRAM) );
  decodeUnit_nbit32 IDU ( .Clk(Clk), .Rst(n1), .en_reg(en_reg_id), .RD1(RD1), 
        .RD2(RD2), .IRAM_instr(IRAM), .PC_Next(PC_Next_fetch), .WR(WR), 
        .ADD_RW(ADD_RW), .DATA_RW(pipe_out), .RW_R_out(RW_R_decode), 
        .RW_I_out(RW_I_decode), .Jump_address(J_imm), .I_immediate_ext_out(
        I_imm), .RD_data_1_out(RD_data_1), .RD_data_2_out(RD_data_2), 
        .PC_Next_out(PC_Next_decode), .Opcode(Opcode), .Func(Func) );
  executionUnit_nbit32 EXE ( .r1(RD_data_1), .r2(RD_data_2), .imm(I_imm), 
        .j_lab(J_imm), .pc(PC_Next_decode), .RW_R(RW_R_decode), .RW_I(
        RW_I_decode), .s2(sel_ex), .s3(sel_mux_rw), .rst(n1), .clk(Clk), 
        .en_reg(en_reg_ex), .alu_sel(alu_sel), .alu_out(alu_out), .r2_out(
        aluR2_to_mem), .b_lab_out(b_from_ex_to_mem), .pc_exe_out(
        pc_from_ex_to_mem), .rw_exe(rw_from_ex_to_mem), .j_lab_out(
        j_from_ex_to_mem) );
  memoryUnit_nbit32 MMU ( .rst(n1), .clk(Clk), .en_reg(en_reg_mem), .b_op(
        b_op_mem), .j_op(j_op_mem), .jal_op(jal_op_mem), .alu_out(alu_out), 
        .r2_out(aluR2_to_mem), .PC(pc_from_ex_to_mem), .lab_b(b_from_ex_to_mem), .lab_j(j_from_ex_to_mem), .rw_exe(rw_from_ex_to_mem), .dataout_from_mem(
        dataout_from_mem), .addr_mem(addr_mem), .datain_mem(datain_mem), 
        .next_PC(pc_from_mem_to_fetch), .alu_out_mem(alu_out_mem), .rw_mem({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, ADD_RW}), .data_out(data_from_mem_to_wb) );
  writeBackUnit_nbit32 WBU ( .MemtoReg(MemtoReg_wb), .ReadData(
        data_from_mem_to_wb), .AluResult(alu_out_mem), .WriteData(pipe_out) );
  BUF_X2 U1 ( .A(Rst), .Z(n1) );
endmodule


module flip_flop_0 ( D, CK, Enable_n, RESET_n, Q );
  input D, CK, Enable_n, RESET_n;
  output Q;
  wire   n1, n4, n2, n3;

  DFFR_X1 Q_reg ( .D(n1), .CK(CK), .RN(RESET_n), .Q(Q), .QN(n4) );
  OAI22_X1 U2 ( .A1(n4), .A2(n3), .B1(Enable_n), .B2(n2), .ZN(n1) );
  INV_X1 U3 ( .A(Enable_n), .ZN(n3) );
  INV_X1 U4 ( .A(D), .ZN(n2) );
endmodule


module flip_flop_1 ( D, CK, Enable_n, RESET_n, Q );
  input D, CK, Enable_n, RESET_n;
  output Q;
  wire   n1, n2, n3, n5;

  DFFR_X1 Q_reg ( .D(n1), .CK(CK), .RN(RESET_n), .Q(Q), .QN(n5) );
  OAI22_X1 U2 ( .A1(n5), .A2(n3), .B1(Enable_n), .B2(n2), .ZN(n1) );
  INV_X1 U3 ( .A(Enable_n), .ZN(n3) );
  INV_X1 U4 ( .A(D), .ZN(n2) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE45_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 ( 
        Clk, Rst, En, IR_opcode, IR_func, PC_OP, EN_REG_IF, EN_REG_ID, RD1, 
        RD2, SEL_EX, EN_REG_EX, SEL_MUX_RW, ALU_OPCODE, EN_REG_MEM, MEM_EN_MEM, 
        RD_MEM, WR_MEM, B_OP_MEM, J_OP_MEM, JAL_OP_MEM, MEM_TO_REG_WB, WR );
  input [5:0] IR_opcode;
  input [10:0] IR_func;
  output [3:0] ALU_OPCODE;
  input Clk, Rst, En;
  output PC_OP, EN_REG_IF, EN_REG_ID, RD1, RD2, SEL_EX, EN_REG_EX, SEL_MUX_RW,
         EN_REG_MEM, MEM_EN_MEM, RD_MEM, WR_MEM, B_OP_MEM, J_OP_MEM,
         JAL_OP_MEM, MEM_TO_REG_WB, WR;
  wire   n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n66, n68, n76, n80,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n65, n67, n69, n70, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103;
  assign PC_OP = 1'b0;
  assign SEL_EX = 1'b0;
  assign SEL_MUX_RW = 1'b0;
  assign RD_MEM = 1'b0;
  assign WR_MEM = 1'b0;
  assign B_OP_MEM = 1'b0;
  assign J_OP_MEM = 1'b0;
  assign JAL_OP_MEM = 1'b0;
  assign WR = 1'b0;

  DFFR_X1 \aluOpcode_3_reg[3]  ( .D(n68), .CK(Clk), .RN(n84), .Q(ALU_OPCODE[3]), .QN(n56) );
  DFFR_X1 \aluOpcode_3_reg[2]  ( .D(n87), .CK(Clk), .RN(n84), .Q(ALU_OPCODE[2]) );
  DFFR_X1 \aluOpcode_3_reg[1]  ( .D(n66), .CK(Clk), .RN(n84), .Q(ALU_OPCODE[1]) );
  DFFR_X1 \aluOpcode_3_reg[0]  ( .D(n80), .CK(Clk), .RN(n84), .Q(ALU_OPCODE[0]), .QN(n76) );
  DFFS_X1 EN_REG_IF_reg ( .D(1'b0), .CK(Clk), .SN(n85), .Q(EN_REG_IF) );
  DFFS_X1 EN_REG_ID_reg ( .D(1'b0), .CK(Clk), .SN(n84), .Q(EN_REG_ID) );
  DFFR_X1 RD1_reg ( .D(1'b1), .CK(Clk), .RN(n84), .Q(RD1) );
  DFFR_X1 RD2_reg ( .D(1'b1), .CK(Clk), .RN(n84), .Q(RD2) );
  DFFS_X1 \cw3_reg[10]  ( .D(n64), .CK(Clk), .SN(n84), .Q(EN_REG_EX), .QN(n55)
         );
  DFFS_X1 \cw3_reg[9]  ( .D(n63), .CK(Clk), .SN(n84), .QN(n53) );
  DFFS_X1 \cw3_reg[2]  ( .D(n62), .CK(Clk), .SN(n85), .QN(n65) );
  DFFS_X1 \cw3_reg[1]  ( .D(n61), .CK(Clk), .SN(n84), .QN(n67) );
  DFFS_X1 \cw4_reg[9]  ( .D(n60), .CK(Clk), .SN(n84), .Q(MEM_EN_MEM), .QN(n54)
         );
  DFFS_X1 \cw4_reg[1]  ( .D(n58), .CK(Clk), .SN(n84), .QN(n69) );
  OAI33_X1 U57 ( .A1(n24), .A2(IR_opcode[1]), .A3(n25), .B1(n26), .B2(n96), 
        .B3(n94), .ZN(n23) );
  XOR2_X1 U58 ( .A(n98), .B(IR_opcode[4]), .Z(n25) );
  OAI33_X1 U59 ( .A1(n88), .A2(IR_func[0]), .A3(n29), .B1(n24), .B2(
        IR_opcode[0]), .B3(n38), .ZN(n37) );
  OAI33_X1 U60 ( .A1(n34), .A2(IR_func[2]), .A3(n103), .B1(n41), .B2(
        IR_opcode[2]), .B3(n98), .ZN(n46) );
  NAND3_X1 U61 ( .A1(n29), .A2(n47), .A3(IR_func[3]), .ZN(n34) );
  NAND3_X1 U71 ( .A1(n89), .A2(n100), .A3(n47), .ZN(n33) );
  NAND3_X1 U72 ( .A1(n97), .A2(n93), .A3(n86), .ZN(n39) );
  NAND3_X1 U73 ( .A1(n86), .A2(IR_opcode[4]), .A3(n52), .ZN(n43) );
  NAND3_X1 U74 ( .A1(n89), .A2(n92), .A3(IR_opcode[2]), .ZN(n24) );
  DFFS_X1 \cw5_reg[1]  ( .D(n57), .CK(Clk), .SN(n85), .Q(MEM_TO_REG_WB), .QN(
        n70) );
  DFFS_X1 \cw4_reg[2]  ( .D(n59), .CK(Clk), .SN(Rst), .Q(EN_REG_MEM), .QN(n83)
         );
  INV_X1 U3 ( .A(n28), .ZN(n88) );
  BUF_X1 U4 ( .A(Rst), .Z(n84) );
  BUF_X1 U5 ( .A(Rst), .Z(n85) );
  NOR2_X1 U6 ( .A1(n101), .A2(n33), .ZN(n28) );
  INV_X1 U7 ( .A(n24), .ZN(n86) );
  INV_X1 U8 ( .A(n34), .ZN(n91) );
  INV_X1 U9 ( .A(n40), .ZN(n96) );
  AND2_X1 U10 ( .A1(n28), .A2(n29), .ZN(n22) );
  INV_X1 U11 ( .A(IR_func[0]), .ZN(n103) );
  INV_X1 U12 ( .A(n27), .ZN(n94) );
  NAND2_X1 U13 ( .A1(n89), .A2(n92), .ZN(n26) );
  INV_X1 U14 ( .A(En), .ZN(n89) );
  NOR4_X1 U15 ( .A1(IR_func[10]), .A2(n96), .A3(n49), .A4(n50), .ZN(n47) );
  OR3_X1 U16 ( .A1(IR_func[7]), .A2(IR_func[6]), .A3(IR_func[4]), .ZN(n49) );
  NAND4_X1 U17 ( .A1(n93), .A2(n92), .A3(n95), .A4(n51), .ZN(n50) );
  NOR3_X1 U18 ( .A1(IR_func[8]), .A2(IR_opcode[1]), .A3(IR_func[9]), .ZN(n51)
         );
  NOR4_X1 U19 ( .A1(IR_func[2]), .A2(n99), .A3(n33), .A4(n102), .ZN(n32) );
  OAI222_X1 U20 ( .A1(En), .A2(n90), .B1(IR_opcode[3]), .B2(n39), .C1(n56), 
        .C2(n89), .ZN(n68) );
  INV_X1 U21 ( .A(n36), .ZN(n90) );
  NOR3_X1 U22 ( .A1(n97), .A2(IR_opcode[4]), .A3(n95), .ZN(n27) );
  OAI22_X1 U23 ( .A1(n40), .A2(n41), .B1(n42), .B2(n34), .ZN(n36) );
  NOR2_X1 U24 ( .A1(IR_func[0]), .A2(IR_func[2]), .ZN(n42) );
  INV_X1 U25 ( .A(IR_func[3]), .ZN(n100) );
  NOR2_X1 U26 ( .A1(n99), .A2(IR_func[1]), .ZN(n29) );
  OAI221_X1 U27 ( .B1(IR_func[0]), .B2(n20), .C1(n76), .C2(n89), .A(n21), .ZN(
        n80) );
  AOI221_X1 U28 ( .B1(n30), .B2(n91), .C1(n31), .C2(n28), .A(n32), .ZN(n20) );
  AOI21_X1 U29 ( .B1(n22), .B2(IR_func[0]), .A(n23), .ZN(n21) );
  NOR2_X1 U30 ( .A1(IR_func[5]), .A2(IR_func[1]), .ZN(n31) );
  NOR2_X1 U31 ( .A1(IR_opcode[2]), .A2(IR_opcode[0]), .ZN(n40) );
  NAND4_X1 U32 ( .A1(n43), .A2(n39), .A3(n44), .A4(n45), .ZN(n66) );
  AOI22_X1 U33 ( .A1(n46), .A2(n89), .B1(En), .B2(ALU_OPCODE[1]), .ZN(n45) );
  OAI21_X1 U34 ( .B1(n48), .B2(n29), .A(n28), .ZN(n44) );
  INV_X1 U35 ( .A(IR_opcode[5]), .ZN(n92) );
  INV_X1 U36 ( .A(IR_opcode[1]), .ZN(n97) );
  INV_X1 U37 ( .A(IR_opcode[3]), .ZN(n95) );
  INV_X1 U38 ( .A(IR_func[2]), .ZN(n101) );
  INV_X1 U39 ( .A(IR_func[5]), .ZN(n99) );
  INV_X1 U40 ( .A(IR_opcode[4]), .ZN(n93) );
  INV_X1 U41 ( .A(n35), .ZN(n87) );
  AOI221_X1 U42 ( .B1(n36), .B2(n89), .C1(En), .C2(ALU_OPCODE[2]), .A(n37), 
        .ZN(n35) );
  AOI21_X1 U43 ( .B1(IR_opcode[4]), .B2(n95), .A(n27), .ZN(n38) );
  NOR3_X1 U44 ( .A1(n102), .A2(IR_func[5]), .A3(IR_func[0]), .ZN(n48) );
  OAI22_X1 U45 ( .A1(n69), .A2(n89), .B1(n67), .B2(En), .ZN(n58) );
  OAI22_X1 U46 ( .A1(n89), .A2(n83), .B1(n65), .B2(En), .ZN(n59) );
  OAI22_X1 U47 ( .A1(n54), .A2(n89), .B1(n53), .B2(En), .ZN(n60) );
  OAI22_X1 U48 ( .A1(n70), .A2(n89), .B1(n69), .B2(En), .ZN(n57) );
  NAND4_X1 U49 ( .A1(IR_opcode[4]), .A2(IR_opcode[3]), .A3(n97), .A4(n92), 
        .ZN(n41) );
  NOR3_X1 U50 ( .A1(n97), .A2(IR_opcode[3]), .A3(IR_opcode[0]), .ZN(n52) );
  NOR2_X1 U51 ( .A1(En), .A2(n101), .ZN(n30) );
  NOR2_X1 U52 ( .A1(n67), .A2(n89), .ZN(n61) );
  NOR2_X1 U53 ( .A1(n65), .A2(n89), .ZN(n62) );
  NOR2_X1 U54 ( .A1(n53), .A2(n89), .ZN(n63) );
  NOR2_X1 U55 ( .A1(n55), .A2(n89), .ZN(n64) );
  INV_X1 U56 ( .A(IR_func[1]), .ZN(n102) );
  INV_X1 U75 ( .A(IR_opcode[0]), .ZN(n98) );
endmodule


module DLX_nbit32 ( Clk, Rst, dout_IRAM, addr_IRAM, MEM_EN_MEM, RD_MEM, WR_MEM, 
        dataout_from_mem, addr_mem, datain_mem, dlx_data_out );
  input [31:0] dout_IRAM;
  output [31:0] addr_IRAM;
  input [31:0] dataout_from_mem;
  output [31:0] addr_mem;
  output [31:0] datain_mem;
  output [31:0] dlx_data_out;
  input Clk, Rst;
  output MEM_EN_MEM, RD_MEM, WR_MEM;
  wire   en_reg_if_i, RD1_i, RD2_i, en_reg_id_i, en_reg_ex_i, en_reg_mem_i,
         MemtoReg_wb_i, CU_en1, CU_en2, n4;
  wire   [5:0] Opcode_i;
  wire   [10:0] Func_i;
  wire   [3:0] alu_sel_i;
  assign RD_MEM = 1'b0;
  assign WR_MEM = 1'b0;

  datapath_nbit32 DataPath_dlx ( .Clk(Clk), .Rst(Rst), .PC_op(1'b0), 
        .en_reg_if(en_reg_if_i), .RD1(RD1_i), .RD2(RD2_i), .dout_IRAM(
        dout_IRAM), .addr_IRAM(addr_IRAM), .en_reg_id(en_reg_id_i), .WR(1'b0), 
        .Opcode(Opcode_i), .Func(Func_i), .sel_ex(1'b0), .sel_mux_rw(1'b0), 
        .en_reg_ex(en_reg_ex_i), .alu_sel(alu_sel_i), .en_reg_mem(en_reg_mem_i), .dataout_from_mem(dataout_from_mem), .addr_mem(addr_mem), .datain_mem(
        datain_mem), .b_op_mem(1'b0), .j_op_mem(1'b0), .jal_op_mem(1'b0), 
        .MemtoReg_wb(MemtoReg_wb_i), .pipe_out(dlx_data_out) );
  flip_flop_0 FF1_en ( .D(n4), .CK(Clk), .Enable_n(1'b0), .RESET_n(1'b1), .Q(
        CU_en1) );
  flip_flop_1 FF2_en ( .D(CU_en1), .CK(Clk), .Enable_n(1'b0), .RESET_n(1'b1), 
        .Q(CU_en2) );
  dlx_cu_MICROCODE_MEM_SIZE45_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 CU_I ( 
        .Clk(Clk), .Rst(Rst), .En(CU_en2), .IR_opcode(Opcode_i), .IR_func(
        Func_i), .EN_REG_IF(en_reg_if_i), .EN_REG_ID(en_reg_id_i), .RD1(RD1_i), 
        .RD2(RD2_i), .EN_REG_EX(en_reg_ex_i), .ALU_OPCODE(alu_sel_i), 
        .EN_REG_MEM(en_reg_mem_i), .MEM_EN_MEM(MEM_EN_MEM), .MEM_TO_REG_WB(
        MemtoReg_wb_i) );
  INV_X1 U14 ( .A(Rst), .ZN(n4) );
endmodule

