
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_nbit32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_nbit32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n14, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U6 : INV_X1 port map( A => n15, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : INV_X1 port map( A => n16, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_1;

architecture SYN_STRUCTURAL of RCA_NBIT4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_2;

architecture SYN_STRUCTURAL of RCA_NBIT4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_4;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n14, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U6 : INV_X1 port map( A => n15, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : INV_X1 port map( A => n16, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_3;

architecture SYN_STRUCTURAL of RCA_NBIT4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_4;

architecture SYN_STRUCTURAL of RCA_NBIT4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_5;

architecture SYN_STRUCTURAL of RCA_NBIT4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_6;

architecture SYN_STRUCTURAL of RCA_NBIT4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_8;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n15, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U6 : INV_X1 port map( A => n14, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_7;

architecture SYN_STRUCTURAL of RCA_NBIT4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_8;

architecture SYN_STRUCTURAL of RCA_NBIT4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_9;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_10;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U6 : INV_X1 port map( A => n17, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U8 : INV_X1 port map( A => n15, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_9;

architecture SYN_STRUCTURAL of RCA_NBIT4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_10;

architecture SYN_STRUCTURAL of RCA_NBIT4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_11;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_12;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n15, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U4 : INV_X1 port map( A => n14, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U6 : INV_X1 port map( A => n17, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U8 : INV_X1 port map( A => n16, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_11;

architecture SYN_STRUCTURAL of RCA_NBIT4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_12;

architecture SYN_STRUCTURAL of RCA_NBIT4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_13;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_14;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n15, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U4 : INV_X1 port map( A => n17, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_13;

architecture SYN_STRUCTURAL of RCA_NBIT4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_14;

architecture SYN_STRUCTURAL of RCA_NBIT4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_15;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => Y(0));
   U2 : INV_X1 port map( A => n15, ZN => Y(1));
   U3 : INV_X1 port map( A => n16, ZN => Y(2));
   U4 : INV_X1 port map( A => n17, ZN => Y(3));
   U5 : INV_X1 port map( A => SEL, ZN => n13);
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_16;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n17, ZN => Y(3));
   U2 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U3 : INV_X1 port map( A => n16, ZN => Y(2));
   U4 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U5 : INV_X1 port map( A => n14, ZN => Y(0));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : INV_X1 port map( A => n15, ZN => Y(1));
   U8 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U9 : INV_X1 port map( A => SEL, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_15;

architecture SYN_STRUCTURAL of RCA_NBIT4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_16;

architecture SYN_STRUCTURAL of RCA_NBIT4_16 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_17;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_18;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_17;

architecture SYN_STRUCTURAL of RCA_NBIT4_17 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_68 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_67 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_66 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_65 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_18;

architecture SYN_STRUCTURAL of RCA_NBIT4_18 is

   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_72 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_71 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_70 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_69 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_19;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_20;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_19;

architecture SYN_STRUCTURAL of RCA_NBIT4_19 is

   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_76 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_75 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_74 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_73 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_20;

architecture SYN_STRUCTURAL of RCA_NBIT4_20 is

   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_80 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_79 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_78 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_77 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_21;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_22;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_21;

architecture SYN_STRUCTURAL of RCA_NBIT4_21 is

   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_84 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_83 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_82 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_81 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_22;

architecture SYN_STRUCTURAL of RCA_NBIT4_22 is

   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_88 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_87 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_86 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_85 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_23;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_24;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n14, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U6 : INV_X1 port map( A => n15, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : INV_X1 port map( A => n16, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_23;

architecture SYN_STRUCTURAL of RCA_NBIT4_23 is

   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_92 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_91 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_90 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_89 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_24;

architecture SYN_STRUCTURAL of RCA_NBIT4_24 is

   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_96 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_95 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_94 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_93 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_25;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_26;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_25;

architecture SYN_STRUCTURAL of RCA_NBIT4_25 is

   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_100 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_99 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_98 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_97 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_26;

architecture SYN_STRUCTURAL of RCA_NBIT4_26 is

   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_104 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_103 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_102 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_101 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_27;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_28;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_27;

architecture SYN_STRUCTURAL of RCA_NBIT4_27 is

   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_108 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_107 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_106 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_105 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_28;

architecture SYN_STRUCTURAL of RCA_NBIT4_28 is

   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_112 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_111 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_110 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_109 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_29;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_30;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_29;

architecture SYN_STRUCTURAL of RCA_NBIT4_29 is

   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_116 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_115 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_114 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_113 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_30;

architecture SYN_STRUCTURAL of RCA_NBIT4_30 is

   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_120 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_119 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_118 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_117 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_31;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => Y(0));
   U2 : INV_X1 port map( A => n15, ZN => Y(1));
   U3 : INV_X1 port map( A => n16, ZN => Y(2));
   U4 : INV_X1 port map( A => n17, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U6 : INV_X1 port map( A => SEL, ZN => n13);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_32;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => Y(0));
   U2 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U5 : INV_X1 port map( A => n16, ZN => Y(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U7 : INV_X1 port map( A => n17, ZN => Y(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U9 : INV_X1 port map( A => SEL, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_31;

architecture SYN_STRUCTURAL of RCA_NBIT4_31 is

   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_124 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_123 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_122 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_121 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_32;

architecture SYN_STRUCTURAL of RCA_NBIT4_32 is

   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_128 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_33;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_34;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_33;

architecture SYN_STRUCTURAL of RCA_NBIT4_33 is

   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_132 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_131 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_130 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_129 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_34;

architecture SYN_STRUCTURAL of RCA_NBIT4_34 is

   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_136 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_135 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_134 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_133 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_35;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_36;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n16, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U4 : INV_X1 port map( A => n17, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U6 : INV_X1 port map( A => n14, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U8 : INV_X1 port map( A => n15, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_35;

architecture SYN_STRUCTURAL of RCA_NBIT4_35 is

   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_140 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_139 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_138 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_137 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_36;

architecture SYN_STRUCTURAL of RCA_NBIT4_36 is

   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_144 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_143 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_142 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_141 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_37;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_38;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_37;

architecture SYN_STRUCTURAL of RCA_NBIT4_37 is

   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_148 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_147 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_146 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_145 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_38;

architecture SYN_STRUCTURAL of RCA_NBIT4_38 is

   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_152 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_151 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_150 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_149 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_39;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_40;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n14, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U6 : INV_X1 port map( A => n15, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : INV_X1 port map( A => n16, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_39;

architecture SYN_STRUCTURAL of RCA_NBIT4_39 is

   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_156 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_155 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_154 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_153 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_40;

architecture SYN_STRUCTURAL of RCA_NBIT4_40 is

   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_160 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_159 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_158 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_157 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_41;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_42;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_41;

architecture SYN_STRUCTURAL of RCA_NBIT4_41 is

   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_164 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_163 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_162 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_161 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_42;

architecture SYN_STRUCTURAL of RCA_NBIT4_42 is

   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_168 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_167 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_166 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_165 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_43;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_44;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_43;

architecture SYN_STRUCTURAL of RCA_NBIT4_43 is

   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_172 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_171 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_170 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_169 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_44;

architecture SYN_STRUCTURAL of RCA_NBIT4_44 is

   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_176 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_175 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_174 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_173 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_45;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_46;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n17, ZN => Y(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_45;

architecture SYN_STRUCTURAL of RCA_NBIT4_45 is

   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_180 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_179 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_178 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_177 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_46;

architecture SYN_STRUCTURAL of RCA_NBIT4_46 is

   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_184 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_183 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_182 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_181 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_47;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => Y(0));
   U2 : INV_X1 port map( A => n15, ZN => Y(1));
   U3 : INV_X1 port map( A => n16, ZN => Y(2));
   U4 : INV_X1 port map( A => n17, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U6 : INV_X1 port map( A => SEL, ZN => n13);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_48;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => Y(0));
   U2 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U5 : INV_X1 port map( A => n16, ZN => Y(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U7 : INV_X1 port map( A => n17, ZN => Y(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U9 : INV_X1 port map( A => SEL, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_47;

architecture SYN_STRUCTURAL of RCA_NBIT4_47 is

   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_188 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_187 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_186 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_185 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_48;

architecture SYN_STRUCTURAL of RCA_NBIT4_48 is

   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_192 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_191 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_190 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_189 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_1;

architecture SYN_structural of CSblock_NBIT4_1 is

   component MUX21_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1000, n_1001, n_1002 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_2 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_1 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1000, Y(2) => 
                           n_1001, Y(1) => n_1002, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_2;

architecture SYN_structural of CSblock_NBIT4_2 is

   component MUX21_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1003, n_1004, n_1005 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_4 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_3 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1003, Y(2) => 
                           n_1004, Y(1) => n_1005, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_3;

architecture SYN_structural of CSblock_NBIT4_3 is

   component MUX21_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1006, n_1007, n_1008 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_6 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_5 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1006, Y(2) => 
                           n_1007, Y(1) => n_1008, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_4;

architecture SYN_structural of CSblock_NBIT4_4 is

   component MUX21_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1009, n_1010, n_1011 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_8 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_7 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1009, Y(2) => 
                           n_1010, Y(1) => n_1011, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_5;

architecture SYN_structural of CSblock_NBIT4_5 is

   component MUX21_GENERIC_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1012, n_1013, n_1014 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_10 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_9 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1012, Y(2) => 
                           n_1013, Y(1) => n_1014, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_6;

architecture SYN_structural of CSblock_NBIT4_6 is

   component MUX21_GENERIC_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1015, n_1016, n_1017 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_12 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_11 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1015, Y(2) => 
                           n_1016, Y(1) => n_1017, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_7;

architecture SYN_structural of CSblock_NBIT4_7 is

   component MUX21_GENERIC_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1018, n_1019, n_1020 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_14 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_13 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1018, Y(2) => 
                           n_1019, Y(1) => n_1020, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_8;

architecture SYN_structural of CSblock_NBIT4_8 is

   component MUX21_GENERIC_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1021, n_1022, n_1023 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_16 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_15 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1021, Y(2) => 
                           n_1022, Y(1) => n_1023, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_1 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_1;

architecture SYN_BEHAVIORAL of GENERAL_G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_2 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_2;

architecture SYN_BEHAVIORAL of GENERAL_G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_3 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_3;

architecture SYN_BEHAVIORAL of GENERAL_G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_4 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_4;

architecture SYN_BEHAVIORAL of GENERAL_G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_1 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_1;

architecture SYN_BEHAVIORAL of GENERAL_PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_2 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_2;

architecture SYN_BEHAVIORAL of GENERAL_PG_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_3 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_3;

architecture SYN_BEHAVIORAL of GENERAL_PG_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_4 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_4;

architecture SYN_BEHAVIORAL of GENERAL_PG_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_5 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_5;

architecture SYN_BEHAVIORAL of GENERAL_G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_6 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_6;

architecture SYN_BEHAVIORAL of GENERAL_G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_5 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_5;

architecture SYN_BEHAVIORAL of GENERAL_PG_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_7 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_7;

architecture SYN_BEHAVIORAL of GENERAL_G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_6 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_6;

architecture SYN_BEHAVIORAL of GENERAL_PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_7 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_7;

architecture SYN_BEHAVIORAL of GENERAL_PG_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_8 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_8;

architecture SYN_BEHAVIORAL of GENERAL_PG_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_9 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_9;

architecture SYN_BEHAVIORAL of GENERAL_PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_10 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_10;

architecture SYN_BEHAVIORAL of GENERAL_PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_11 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_11;

architecture SYN_BEHAVIORAL of GENERAL_PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_12 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_12;

architecture SYN_BEHAVIORAL of GENERAL_PG_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_13 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_13;

architecture SYN_BEHAVIORAL of GENERAL_PG_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_14 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_14;

architecture SYN_BEHAVIORAL of GENERAL_PG_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_15 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_15;

architecture SYN_BEHAVIORAL of GENERAL_PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_16 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_16;

architecture SYN_BEHAVIORAL of GENERAL_PG_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_17 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_17;

architecture SYN_BEHAVIORAL of GENERAL_PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_18 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_18;

architecture SYN_BEHAVIORAL of GENERAL_PG_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_19 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_19;

architecture SYN_BEHAVIORAL of GENERAL_PG_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_20 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_20;

architecture SYN_BEHAVIORAL of GENERAL_PG_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_21 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_21;

architecture SYN_BEHAVIORAL of GENERAL_PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_22 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_22;

architecture SYN_BEHAVIORAL of GENERAL_PG_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_23 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_23;

architecture SYN_BEHAVIORAL of GENERAL_PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_24 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_24;

architecture SYN_BEHAVIORAL of GENERAL_PG_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_25 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_25;

architecture SYN_BEHAVIORAL of GENERAL_PG_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_26 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_26;

architecture SYN_BEHAVIORAL of GENERAL_PG_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_8 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_8;

architecture SYN_BEHAVIORAL of GENERAL_G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_27 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_27;

architecture SYN_BEHAVIORAL of GENERAL_PG_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_9 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_9;

architecture SYN_BEHAVIORAL of GENERAL_G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_1 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_1;

architecture SYN_BEHAVIORAL of PG_block_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_2 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_2;

architecture SYN_BEHAVIORAL of PG_block_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_3 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_3;

architecture SYN_BEHAVIORAL of PG_block_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_4 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_4;

architecture SYN_BEHAVIORAL of PG_block_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_5 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_5;

architecture SYN_BEHAVIORAL of PG_block_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_6 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_6;

architecture SYN_BEHAVIORAL of PG_block_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_7 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_7;

architecture SYN_BEHAVIORAL of PG_block_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_8 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_8;

architecture SYN_BEHAVIORAL of PG_block_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_9 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_9;

architecture SYN_BEHAVIORAL of PG_block_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_10 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_10;

architecture SYN_BEHAVIORAL of PG_block_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_11 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_11;

architecture SYN_BEHAVIORAL of PG_block_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_12 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_12;

architecture SYN_BEHAVIORAL of PG_block_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_13 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_13;

architecture SYN_BEHAVIORAL of PG_block_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_14 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_14;

architecture SYN_BEHAVIORAL of PG_block_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_15 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_15;

architecture SYN_BEHAVIORAL of PG_block_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_16 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_16;

architecture SYN_BEHAVIORAL of PG_block_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_17 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_17;

architecture SYN_BEHAVIORAL of PG_block_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_18 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_18;

architecture SYN_BEHAVIORAL of PG_block_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_19 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_19;

architecture SYN_BEHAVIORAL of PG_block_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_20 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_20;

architecture SYN_BEHAVIORAL of PG_block_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_21 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_21;

architecture SYN_BEHAVIORAL of PG_block_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_22 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_22;

architecture SYN_BEHAVIORAL of PG_block_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_23 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_23;

architecture SYN_BEHAVIORAL of PG_block_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_24 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_24;

architecture SYN_BEHAVIORAL of PG_block_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_25 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_25;

architecture SYN_BEHAVIORAL of PG_block_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_26 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_26;

architecture SYN_BEHAVIORAL of PG_block_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_27 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_27;

architecture SYN_BEHAVIORAL of PG_block_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_28 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_28;

architecture SYN_BEHAVIORAL of PG_block_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_29 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_29;

architecture SYN_BEHAVIORAL of PG_block_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_30 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_30;

architecture SYN_BEHAVIORAL of PG_block_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_31 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_31;

architecture SYN_BEHAVIORAL of PG_block_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_10 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_10;

architecture SYN_BEHAVIORAL of GENERAL_G_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_32 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_32;

architecture SYN_BEHAVIORAL of PG_block_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_49;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_50;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_49;

architecture SYN_STRUCTURAL of RCA_NBIT4_49 is

   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_196 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_195 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_194 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_193 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_50;

architecture SYN_STRUCTURAL of RCA_NBIT4_50 is

   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_200 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_199 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_198 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_197 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_51;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_52;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_51;

architecture SYN_STRUCTURAL of RCA_NBIT4_51 is

   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_204 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_203 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_202 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_201 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_52;

architecture SYN_STRUCTURAL of RCA_NBIT4_52 is

   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_208 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_207 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_206 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_205 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_53;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_54;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_53;

architecture SYN_STRUCTURAL of RCA_NBIT4_53 is

   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_212 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_211 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_210 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_209 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_54;

architecture SYN_STRUCTURAL of RCA_NBIT4_54 is

   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_216 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_215 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_214 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_213 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_55;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_56;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n15, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U6 : INV_X1 port map( A => n17, ZN => Y(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_55;

architecture SYN_STRUCTURAL of RCA_NBIT4_55 is

   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_220 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_219 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_218 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_217 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_56;

architecture SYN_STRUCTURAL of RCA_NBIT4_56 is

   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_224 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_223 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_222 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_221 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_57;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_58;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_57;

architecture SYN_STRUCTURAL of RCA_NBIT4_57 is

   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_228 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_227 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_226 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_225 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_58;

architecture SYN_STRUCTURAL of RCA_NBIT4_58 is

   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_232 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_231 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_230 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_229 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_59;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_60;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_59;

architecture SYN_STRUCTURAL of RCA_NBIT4_59 is

   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_236 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_235 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_234 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_233 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_60;

architecture SYN_STRUCTURAL of RCA_NBIT4_60 is

   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_240 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_239 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_238 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_237 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_61;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n14, ZN => Y(0));
   U3 : INV_X1 port map( A => n15, ZN => Y(1));
   U4 : INV_X1 port map( A => n16, ZN => Y(2));
   U5 : INV_X1 port map( A => n17, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_62;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n13);
   U2 : INV_X1 port map( A => n17, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n17);
   U4 : INV_X1 port map( A => n15, ZN => Y(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n15);
   U6 : INV_X1 port map( A => n16, ZN => Y(2));
   U7 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n16);
   U8 : INV_X1 port map( A => n14, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_61;

architecture SYN_STRUCTURAL of RCA_NBIT4_61 is

   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_244 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_243 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_242 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_241 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_62;

architecture SYN_STRUCTURAL of RCA_NBIT4_62 is

   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_248 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_247 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_246 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_245 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_63;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => Y(0));
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : INV_X1 port map( A => n7, ZN => Y(2));
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U6 : INV_X1 port map( A => SEL, ZN => n13);
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U8 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => Y(0));
   U2 : AOI22_X1 port map( A1 => A(0), A2 => n13, B1 => B(0), B2 => SEL, ZN => 
                           n9);
   U3 : INV_X1 port map( A => n8, ZN => Y(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n13, B1 => B(1), B2 => SEL, ZN => 
                           n8);
   U5 : INV_X1 port map( A => n7, ZN => Y(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n13, B1 => B(2), B2 => SEL, ZN => 
                           n7);
   U7 : INV_X1 port map( A => n6, ZN => Y(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n13, B1 => SEL, B2 => B(3), ZN => 
                           n6);
   U9 : INV_X1 port map( A => SEL, ZN => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_63;

architecture SYN_STRUCTURAL of RCA_NBIT4_63 is

   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_252 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_251 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_250 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_249 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity RCA_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_0;

architecture SYN_STRUCTURAL of RCA_NBIT4_0 is

   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_255 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_254 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_253 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_9;

architecture SYN_structural of CSblock_NBIT4_9 is

   component MUX21_GENERIC_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1024, n_1025, n_1026 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_18 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_17 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1024, Y(2) => 
                           n_1025, Y(1) => n_1026, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_10;

architecture SYN_structural of CSblock_NBIT4_10 is

   component MUX21_GENERIC_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1027, n_1028, n_1029 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_20 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_19 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1027, Y(2) => 
                           n_1028, Y(1) => n_1029, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_11;

architecture SYN_structural of CSblock_NBIT4_11 is

   component MUX21_GENERIC_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1030, n_1031, n_1032 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_22 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_21 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1030, Y(2) => 
                           n_1031, Y(1) => n_1032, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_12;

architecture SYN_structural of CSblock_NBIT4_12 is

   component MUX21_GENERIC_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1033, n_1034, n_1035 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_24 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_23 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1033, Y(2) => 
                           n_1034, Y(1) => n_1035, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_13;

architecture SYN_structural of CSblock_NBIT4_13 is

   component MUX21_GENERIC_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1036, n_1037, n_1038 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_26 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_25 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1036, Y(2) => 
                           n_1037, Y(1) => n_1038, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_14;

architecture SYN_structural of CSblock_NBIT4_14 is

   component MUX21_GENERIC_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1039, n_1040, n_1041 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_28 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_27 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1039, Y(2) => 
                           n_1040, Y(1) => n_1041, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_15;

architecture SYN_structural of CSblock_NBIT4_15 is

   component MUX21_GENERIC_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1042, n_1043, n_1044 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_30 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_29 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1042, Y(2) => 
                           n_1043, Y(1) => n_1044, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_16;

architecture SYN_structural of CSblock_NBIT4_16 is

   component MUX21_GENERIC_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1045, n_1046, n_1047 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_31 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_32 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_31 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1045, Y(2) => 
                           n_1046, Y(1) => n_1047, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_11 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_11;

architecture SYN_BEHAVIORAL of GENERAL_G_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_12 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_12;

architecture SYN_BEHAVIORAL of GENERAL_G_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_13 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_13;

architecture SYN_BEHAVIORAL of GENERAL_G_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_14 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_14;

architecture SYN_BEHAVIORAL of GENERAL_G_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_28 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_28;

architecture SYN_BEHAVIORAL of GENERAL_PG_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_29 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_29;

architecture SYN_BEHAVIORAL of GENERAL_PG_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_30 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_30;

architecture SYN_BEHAVIORAL of GENERAL_PG_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_31 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_31;

architecture SYN_BEHAVIORAL of GENERAL_PG_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_15 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_15;

architecture SYN_BEHAVIORAL of GENERAL_G_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_16 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_16;

architecture SYN_BEHAVIORAL of GENERAL_G_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_32 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_32;

architecture SYN_BEHAVIORAL of GENERAL_PG_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_17 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_17;

architecture SYN_BEHAVIORAL of GENERAL_G_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_33 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_33;

architecture SYN_BEHAVIORAL of GENERAL_PG_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_34 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_34;

architecture SYN_BEHAVIORAL of GENERAL_PG_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_35 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_35;

architecture SYN_BEHAVIORAL of GENERAL_PG_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_36 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_36;

architecture SYN_BEHAVIORAL of GENERAL_PG_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_37 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_37;

architecture SYN_BEHAVIORAL of GENERAL_PG_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_38 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_38;

architecture SYN_BEHAVIORAL of GENERAL_PG_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_39 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_39;

architecture SYN_BEHAVIORAL of GENERAL_PG_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_40 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_40;

architecture SYN_BEHAVIORAL of GENERAL_PG_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_41 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_41;

architecture SYN_BEHAVIORAL of GENERAL_PG_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_42 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_42;

architecture SYN_BEHAVIORAL of GENERAL_PG_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_43 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_43;

architecture SYN_BEHAVIORAL of GENERAL_PG_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_44 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_44;

architecture SYN_BEHAVIORAL of GENERAL_PG_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_45 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_45;

architecture SYN_BEHAVIORAL of GENERAL_PG_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_46 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_46;

architecture SYN_BEHAVIORAL of GENERAL_PG_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_47 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_47;

architecture SYN_BEHAVIORAL of GENERAL_PG_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_48 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_48;

architecture SYN_BEHAVIORAL of GENERAL_PG_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_49 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_49;

architecture SYN_BEHAVIORAL of GENERAL_PG_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_50 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_50;

architecture SYN_BEHAVIORAL of GENERAL_PG_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_51 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_51;

architecture SYN_BEHAVIORAL of GENERAL_PG_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_52 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_52;

architecture SYN_BEHAVIORAL of GENERAL_PG_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_53 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_53;

architecture SYN_BEHAVIORAL of GENERAL_PG_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_18 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_18;

architecture SYN_BEHAVIORAL of GENERAL_G_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_54 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_54;

architecture SYN_BEHAVIORAL of GENERAL_PG_54 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_19 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_19;

architecture SYN_BEHAVIORAL of GENERAL_G_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_33 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_33;

architecture SYN_BEHAVIORAL of PG_block_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_34 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_34;

architecture SYN_BEHAVIORAL of PG_block_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_35 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_35;

architecture SYN_BEHAVIORAL of PG_block_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_36 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_36;

architecture SYN_BEHAVIORAL of PG_block_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_37 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_37;

architecture SYN_BEHAVIORAL of PG_block_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_38 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_38;

architecture SYN_BEHAVIORAL of PG_block_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_39 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_39;

architecture SYN_BEHAVIORAL of PG_block_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_40 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_40;

architecture SYN_BEHAVIORAL of PG_block_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_41 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_41;

architecture SYN_BEHAVIORAL of PG_block_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_42 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_42;

architecture SYN_BEHAVIORAL of PG_block_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_43 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_43;

architecture SYN_BEHAVIORAL of PG_block_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_44 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_44;

architecture SYN_BEHAVIORAL of PG_block_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_45 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_45;

architecture SYN_BEHAVIORAL of PG_block_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_46 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_46;

architecture SYN_BEHAVIORAL of PG_block_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_47 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_47;

architecture SYN_BEHAVIORAL of PG_block_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_48 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_48;

architecture SYN_BEHAVIORAL of PG_block_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_49 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_49;

architecture SYN_BEHAVIORAL of PG_block_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_50 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_50;

architecture SYN_BEHAVIORAL of PG_block_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_51 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_51;

architecture SYN_BEHAVIORAL of PG_block_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_52 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_52;

architecture SYN_BEHAVIORAL of PG_block_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_53 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_53;

architecture SYN_BEHAVIORAL of PG_block_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_54 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_54;

architecture SYN_BEHAVIORAL of PG_block_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_55 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_55;

architecture SYN_BEHAVIORAL of PG_block_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_56 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_56;

architecture SYN_BEHAVIORAL of PG_block_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_57 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_57;

architecture SYN_BEHAVIORAL of PG_block_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_58 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_58;

architecture SYN_BEHAVIORAL of PG_block_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_59 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_59;

architecture SYN_BEHAVIORAL of PG_block_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_60 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_60;

architecture SYN_BEHAVIORAL of PG_block_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_61 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_61;

architecture SYN_BEHAVIORAL of PG_block_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_62 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_62;

architecture SYN_BEHAVIORAL of PG_block_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_63 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_63;

architecture SYN_BEHAVIORAL of PG_block_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_20 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_20;

architecture SYN_BEHAVIORAL of GENERAL_G_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_64 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_64;

architecture SYN_BEHAVIORAL of PG_block_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_17;

architecture SYN_structural of CSblock_NBIT4_17 is

   component MUX21_GENERIC_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1048, n_1049, n_1050 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_34 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_33 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_34 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_33 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1048, Y(2) => 
                           n_1049, Y(1) => n_1050, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_18;

architecture SYN_structural of CSblock_NBIT4_18 is

   component MUX21_GENERIC_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1051, n_1052, n_1053 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_36 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_35 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_36 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_35 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1051, Y(2) => 
                           n_1052, Y(1) => n_1053, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_19;

architecture SYN_structural of CSblock_NBIT4_19 is

   component MUX21_GENERIC_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1054, n_1055, n_1056 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_38 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_37 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_38 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_37 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1054, Y(2) => 
                           n_1055, Y(1) => n_1056, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_20;

architecture SYN_structural of CSblock_NBIT4_20 is

   component MUX21_GENERIC_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1057, n_1058, n_1059 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_39 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_40 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_39 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1057, Y(2) => 
                           n_1058, Y(1) => n_1059, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_21;

architecture SYN_structural of CSblock_NBIT4_21 is

   component MUX21_GENERIC_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1060, n_1061, n_1062 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_42 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_41 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_42 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_41 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1060, Y(2) => 
                           n_1061, Y(1) => n_1062, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_22;

architecture SYN_structural of CSblock_NBIT4_22 is

   component MUX21_GENERIC_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1063, n_1064, n_1065 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_44 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_43 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_44 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_43 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1063, Y(2) => 
                           n_1064, Y(1) => n_1065, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_23;

architecture SYN_structural of CSblock_NBIT4_23 is

   component MUX21_GENERIC_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1066, n_1067, n_1068 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_46 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_45 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_46 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_45 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1066, Y(2) => 
                           n_1067, Y(1) => n_1068, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_24;

architecture SYN_structural of CSblock_NBIT4_24 is

   component MUX21_GENERIC_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1069, n_1070, n_1071 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_47 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_48 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_47 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1069, Y(2) => 
                           n_1070, Y(1) => n_1071, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_21 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_21;

architecture SYN_BEHAVIORAL of GENERAL_G_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_22 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_22;

architecture SYN_BEHAVIORAL of GENERAL_G_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_23 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_23;

architecture SYN_BEHAVIORAL of GENERAL_G_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_24 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_24;

architecture SYN_BEHAVIORAL of GENERAL_G_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_55 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_55;

architecture SYN_BEHAVIORAL of GENERAL_PG_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_56 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_56;

architecture SYN_BEHAVIORAL of GENERAL_PG_56 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_57 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_57;

architecture SYN_BEHAVIORAL of GENERAL_PG_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_58 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_58;

architecture SYN_BEHAVIORAL of GENERAL_PG_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_25 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_25;

architecture SYN_BEHAVIORAL of GENERAL_G_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_26 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_26;

architecture SYN_BEHAVIORAL of GENERAL_G_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_59 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_59;

architecture SYN_BEHAVIORAL of GENERAL_PG_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_27 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_27;

architecture SYN_BEHAVIORAL of GENERAL_G_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_60 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_60;

architecture SYN_BEHAVIORAL of GENERAL_PG_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_61 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_61;

architecture SYN_BEHAVIORAL of GENERAL_PG_61 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_62 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_62;

architecture SYN_BEHAVIORAL of GENERAL_PG_62 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_63 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_63;

architecture SYN_BEHAVIORAL of GENERAL_PG_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_64 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_64;

architecture SYN_BEHAVIORAL of GENERAL_PG_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_65 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_65;

architecture SYN_BEHAVIORAL of GENERAL_PG_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_66 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_66;

architecture SYN_BEHAVIORAL of GENERAL_PG_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_67 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_67;

architecture SYN_BEHAVIORAL of GENERAL_PG_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_68 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_68;

architecture SYN_BEHAVIORAL of GENERAL_PG_68 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_69 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_69;

architecture SYN_BEHAVIORAL of GENERAL_PG_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_70 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_70;

architecture SYN_BEHAVIORAL of GENERAL_PG_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_71 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_71;

architecture SYN_BEHAVIORAL of GENERAL_PG_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_72 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_72;

architecture SYN_BEHAVIORAL of GENERAL_PG_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_73 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_73;

architecture SYN_BEHAVIORAL of GENERAL_PG_73 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_74 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_74;

architecture SYN_BEHAVIORAL of GENERAL_PG_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_75 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_75;

architecture SYN_BEHAVIORAL of GENERAL_PG_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_76 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_76;

architecture SYN_BEHAVIORAL of GENERAL_PG_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_77 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_77;

architecture SYN_BEHAVIORAL of GENERAL_PG_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_78 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_78;

architecture SYN_BEHAVIORAL of GENERAL_PG_78 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_79 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_79;

architecture SYN_BEHAVIORAL of GENERAL_PG_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_80 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_80;

architecture SYN_BEHAVIORAL of GENERAL_PG_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_28 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_28;

architecture SYN_BEHAVIORAL of GENERAL_G_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_81 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_81;

architecture SYN_BEHAVIORAL of GENERAL_PG_81 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_29 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_29;

architecture SYN_BEHAVIORAL of GENERAL_G_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_65 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_65;

architecture SYN_BEHAVIORAL of PG_block_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_66 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_66;

architecture SYN_BEHAVIORAL of PG_block_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_67 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_67;

architecture SYN_BEHAVIORAL of PG_block_67 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_68 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_68;

architecture SYN_BEHAVIORAL of PG_block_68 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_69 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_69;

architecture SYN_BEHAVIORAL of PG_block_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_70 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_70;

architecture SYN_BEHAVIORAL of PG_block_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_71 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_71;

architecture SYN_BEHAVIORAL of PG_block_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_72 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_72;

architecture SYN_BEHAVIORAL of PG_block_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_73 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_73;

architecture SYN_BEHAVIORAL of PG_block_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_74 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_74;

architecture SYN_BEHAVIORAL of PG_block_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_75 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_75;

architecture SYN_BEHAVIORAL of PG_block_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_76 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_76;

architecture SYN_BEHAVIORAL of PG_block_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_77 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_77;

architecture SYN_BEHAVIORAL of PG_block_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_78 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_78;

architecture SYN_BEHAVIORAL of PG_block_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_79 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_79;

architecture SYN_BEHAVIORAL of PG_block_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_80 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_80;

architecture SYN_BEHAVIORAL of PG_block_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_81 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_81;

architecture SYN_BEHAVIORAL of PG_block_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_82 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_82;

architecture SYN_BEHAVIORAL of PG_block_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_83 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_83;

architecture SYN_BEHAVIORAL of PG_block_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_84 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_84;

architecture SYN_BEHAVIORAL of PG_block_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_85 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_85;

architecture SYN_BEHAVIORAL of PG_block_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_86 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_86;

architecture SYN_BEHAVIORAL of PG_block_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_87 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_87;

architecture SYN_BEHAVIORAL of PG_block_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_88 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_88;

architecture SYN_BEHAVIORAL of PG_block_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_89 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_89;

architecture SYN_BEHAVIORAL of PG_block_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_90 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_90;

architecture SYN_BEHAVIORAL of PG_block_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_91 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_91;

architecture SYN_BEHAVIORAL of PG_block_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_92 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_92;

architecture SYN_BEHAVIORAL of PG_block_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_93 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_93;

architecture SYN_BEHAVIORAL of PG_block_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_94 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_94;

architecture SYN_BEHAVIORAL of PG_block_94 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_95 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_95;

architecture SYN_BEHAVIORAL of PG_block_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_30 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_30;

architecture SYN_BEHAVIORAL of GENERAL_G_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_96 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_96;

architecture SYN_BEHAVIORAL of PG_block_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity comparator_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_DW01_cmp6_0;

architecture SYN_rpl of comparator_DW01_cmp6_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n202, n292, n65, n66, n69, n71, n72, n74, n75, n77, n80, n81, n83, 
      n84, n86, n87, n89, n92, n93, n95, n96, n98, n99, n101, n104, n105, n108,
      n110, n111, n113, n116, n117, n120, n122, n123, n125, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      net52631, net52642, net52646, net52650, net52651, net52652, net54692, 
      n203, n204, n205, n206, n207, n208, n209, n210, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291 : std_logic;

begin
   
   U101 : XOR2_X1 port map( A => A(30), B => net52651, Z => n69);
   U170 : NAND3_X1 port map( A1 => n196, A2 => n149, A3 => n146, ZN => n195);
   U174 : NAND3_X1 port map( A1 => n199, A2 => n198, A3 => n283, ZN => n196);
   U1 : AND2_X1 port map( A1 => n89, A2 => n92, ZN => n226);
   U2 : NAND2_X1 port map( A1 => n86, A2 => n207, ZN => n228);
   U3 : NOR2_X1 port map( A1 => n84, A2 => n81, ZN => n244);
   U4 : NAND2_X1 port map( A1 => n83, A2 => n243, ZN => n242);
   U5 : INV_X1 port map( A => n87, ZN => n243);
   U6 : NAND2_X1 port map( A1 => n125, A2 => n128, ZN => n216);
   U7 : OAI21_X1 port map( B1 => n215, B2 => n234, A => n235, ZN => n219);
   U8 : NOR2_X1 port map( A1 => n123, A2 => n208, ZN => n235);
   U9 : NAND2_X1 port map( A1 => n122, A2 => n203, ZN => n234);
   U10 : NOR2_X1 port map( A1 => n210, A2 => n216, ZN => n215);
   U11 : NOR2_X1 port map( A1 => n120, A2 => n117, ZN => n218);
   U12 : NAND2_X1 port map( A1 => n113, A2 => n116, ZN => n220);
   U13 : OAI21_X1 port map( B1 => n217, B2 => n236, A => n237, ZN => n248);
   U14 : NOR2_X1 port map( A1 => n111, A2 => n209, ZN => n237);
   U15 : NAND2_X1 port map( A1 => n110, A2 => n205, ZN => n236);
   U16 : AOI21_X1 port map( B1 => n218, B2 => n219, A => n220, ZN => n217);
   U17 : NOR2_X1 port map( A1 => n108, A2 => n105, ZN => n238);
   U18 : AOI21_X1 port map( B1 => n222, B2 => n223, A => n224, ZN => n221);
   U19 : AND2_X1 port map( A1 => n101, A2 => n104, ZN => n222);
   U20 : NAND2_X1 port map( A1 => n98, A2 => n206, ZN => n224);
   U21 : NAND2_X1 port map( A1 => n238, A2 => n248, ZN => n223);
   U22 : NOR2_X1 port map( A1 => n96, A2 => n93, ZN => n241);
   U23 : NAND2_X1 port map( A1 => n95, A2 => n240, ZN => n239);
   U24 : INV_X1 port map( A => n99, ZN => n240);
   U25 : AND2_X1 port map( A1 => n77, A2 => n80, ZN => n230);
   U26 : NAND2_X1 port map( A1 => n74, A2 => n204, ZN => n232);
   U27 : NOR2_X1 port map( A1 => n72, A2 => n233, ZN => n247);
   U28 : INV_X1 port map( A => n69, ZN => n233);
   U29 : NAND2_X1 port map( A1 => n71, A2 => n246, ZN => n245);
   U30 : INV_X1 port map( A => n75, ZN => n246);
   U31 : OR2_X1 port map( A1 => n262, A2 => B(11), ZN => n203);
   U32 : OR2_X1 port map( A1 => n273, A2 => B(27), ZN => n204);
   U33 : OR2_X1 port map( A1 => n289, A2 => B(15), ZN => n205);
   U34 : OR2_X1 port map( A1 => n287, A2 => B(19), ZN => n206);
   U35 : OR2_X1 port map( A1 => n269, A2 => B(23), ZN => n207);
   U36 : AND2_X1 port map( A1 => B(13), A2 => n263, ZN => n208);
   U37 : AND2_X1 port map( A1 => B(17), A2 => n265, ZN => n209);
   U38 : AND2_X1 port map( A1 => n127, A2 => net52631, ZN => n210);
   U39 : CLKBUF_X1 port map( A => n276, Z => LE);
   U40 : AOI21_X1 port map( B1 => n230, B2 => n231, A => n232, ZN => n229);
   U41 : OAI21_X1 port map( B1 => n225, B2 => n242, A => n244, ZN => n231);
   U42 : NAND2_X1 port map( A1 => n213, A2 => n214, ZN => net52652);
   U43 : AOI21_X1 port map( B1 => n226, B2 => n227, A => n228, ZN => n225);
   U44 : NOR2_X1 port map( A1 => n252, A2 => B(0), ZN => n212);
   U45 : OAI21_X1 port map( B1 => n229, B2 => n245, A => n247, ZN => n214);
   U46 : OAI21_X1 port map( B1 => n221, B2 => n239, A => n241, ZN => n227);
   U47 : NAND2_X1 port map( A1 => B(30), A2 => net54692, ZN => n213);
   U48 : OR2_X1 port map( A1 => B(2), A2 => n253, ZN => n198);
   U49 : AOI21_X1 port map( B1 => net52652, B2 => n65, A => n66, ZN => GE);
   U50 : NAND2_X1 port map( A1 => B(0), A2 => n250, ZN => n154);
   U51 : AND2_X1 port map( A1 => n252, A2 => n251, ZN => n250);
   U52 : INV_X1 port map( A => A(1), ZN => n251);
   U53 : NOR2_X1 port map( A1 => n192, A2 => n135, ZN => n134);
   U54 : NOR2_X1 port map( A1 => n192, A2 => n132, ZN => n188);
   U55 : INV_X1 port map( A => n95, ZN => net52642);
   U56 : INV_X1 port map( A => n131, ZN => n278);
   U57 : INV_X1 port map( A => n141, ZN => n281);
   U58 : INV_X1 port map( A => n129, ZN => net52631);
   U59 : OAI211_X1 port map( C1 => n166, C2 => n167, A => n89, B => n86, ZN => 
                           n165);
   U60 : NAND2_X1 port map( A1 => n207, A2 => n169, ZN => n167);
   U61 : AOI211_X1 port map( C1 => n171, C2 => n170, A => n93, B => net52642, 
                           ZN => n166);
   U62 : OAI211_X1 port map( C1 => n160, C2 => n161, A => n77, B => n74, ZN => 
                           n159);
   U63 : NAND2_X1 port map( A1 => n204, A2 => n163, ZN => n161);
   U64 : AOI211_X1 port map( C1 => n165, C2 => n164, A => n81, B => net52646, 
                           ZN => n160);
   U65 : OAI211_X1 port map( C1 => n178, C2 => n179, A => n113, B => n110, ZN 
                           => n177);
   U66 : NAND2_X1 port map( A1 => n205, A2 => n181, ZN => n179);
   U67 : AOI211_X1 port map( C1 => n183, C2 => n182, A => n117, B => n208, ZN 
                           => n178);
   U68 : OAI211_X1 port map( C1 => n184, C2 => n185, A => n125, B => n122, ZN 
                           => n183);
   U69 : NAND2_X1 port map( A1 => n203, A2 => n187, ZN => n185);
   U70 : AOI211_X1 port map( C1 => n189, C2 => n188, A => n129, B => n278, ZN 
                           => n184);
   U71 : NOR2_X1 port map( A1 => n260, A2 => B(9), ZN => n132);
   U72 : OAI211_X1 port map( C1 => n172, C2 => n173, A => n101, B => n98, ZN =>
                           n171);
   U73 : NAND2_X1 port map( A1 => n206, A2 => n175, ZN => n173);
   U74 : AOI211_X1 port map( C1 => n177, C2 => n176, A => n105, B => n209, ZN 
                           => n172);
   U75 : NOR2_X1 port map( A1 => n162, A2 => n75, ZN => n74);
   U76 : NOR2_X1 port map( A1 => n186, A2 => n123, ZN => n122);
   U77 : NOR2_X1 port map( A1 => n180, A2 => n111, ZN => n110);
   U78 : NOR2_X1 port map( A1 => n174, A2 => n99, ZN => n98);
   U79 : NOR2_X1 port map( A1 => n168, A2 => n87, ZN => n86);
   U80 : NAND2_X1 port map( A1 => B(9), A2 => n260, ZN => n131);
   U81 : NOR2_X1 port map( A1 => n197, A2 => n147, ZN => n146);
   U82 : NOR2_X1 port map( A1 => n162, A2 => n72, ZN => n158);
   U83 : NOR2_X1 port map( A1 => n197, A2 => n144, ZN => n194);
   U84 : NOR2_X1 port map( A1 => n186, A2 => n120, ZN => n182);
   U85 : NOR2_X1 port map( A1 => n180, A2 => n108, ZN => n176);
   U86 : NOR2_X1 port map( A1 => n174, A2 => n96, ZN => n170);
   U87 : NOR2_X1 port map( A1 => n168, A2 => n84, ZN => n164);
   U88 : NAND2_X1 port map( A1 => n169, A2 => n92, ZN => n93);
   U89 : NAND2_X1 port map( A1 => n163, A2 => n80, ZN => n81);
   U90 : NAND2_X1 port map( A1 => n193, A2 => n140, ZN => n141);
   U91 : NAND2_X1 port map( A1 => n187, A2 => n128, ZN => n129);
   U92 : NAND2_X1 port map( A1 => n175, A2 => n104, ZN => n105);
   U93 : NAND2_X1 port map( A1 => n181, A2 => n116, ZN => n117);
   U94 : AND2_X1 port map( A1 => n198, A2 => n153, ZN => n152);
   U95 : INV_X1 port map( A => n143, ZN => n282);
   U96 : INV_X1 port map( A => n83, ZN => net52646);
   U97 : INV_X1 port map( A => n140, ZN => n280);
   U98 : INV_X1 port map( A => n153, ZN => n284);
   U99 : NOR2_X1 port map( A1 => n255, A2 => B(4), ZN => n197);
   U100 : NOR2_X1 port map( A1 => n288, A2 => B(16), ZN => n180);
   U102 : NOR2_X1 port map( A1 => n270, A2 => B(24), ZN => n168);
   U103 : NOR2_X1 port map( A1 => n291, A2 => B(12), ZN => n186);
   U104 : NOR2_X1 port map( A1 => n290, A2 => B(20), ZN => n174);
   U105 : NOR2_X1 port map( A1 => n275, A2 => B(29), ZN => n72);
   U106 : NOR2_X1 port map( A1 => n254, A2 => B(3), ZN => n150);
   U107 : OAI211_X1 port map( C1 => n190, C2 => n191, A => n137, B => n134, ZN 
                           => n189);
   U108 : NAND2_X1 port map( A1 => n279, A2 => n193, ZN => n191);
   U109 : AOI211_X1 port map( C1 => n194, C2 => n195, A => n141, B => n282, ZN 
                           => n190);
   U110 : INV_X1 port map( A => n138, ZN => n279);
   U111 : NOR2_X1 port map( A1 => n256, A2 => B(5), ZN => n144);
   U112 : NAND2_X1 port map( A1 => B(3), A2 => n254, ZN => n149);
   U113 : NOR2_X1 port map( A1 => n258, A2 => B(7), ZN => n138);
   U114 : NOR2_X1 port map( A1 => n265, A2 => B(17), ZN => n108);
   U115 : NOR2_X1 port map( A1 => n271, A2 => B(25), ZN => n84);
   U116 : NAND2_X1 port map( A1 => B(6), A2 => n257, ZN => n140);
   U117 : NAND2_X1 port map( A1 => B(26), A2 => n272, ZN => n80);
   U118 : NAND2_X1 port map( A1 => B(19), A2 => n287, ZN => n101);
   U119 : NAND2_X1 port map( A1 => B(29), A2 => n275, ZN => n71);
   U120 : OAI21_X1 port map( B1 => n156, B2 => n66, A => n65, ZN => n202);
   U121 : AOI22_X1 port map( A1 => A(30), A2 => net52651, B1 => n157, B2 => n69
                           , ZN => n156);
   U122 : AOI21_X1 port map( B1 => n159, B2 => n158, A => net52650, ZN => n157)
                           ;
   U123 : INV_X1 port map( A => n71, ZN => net52650);
   U124 : NAND2_X1 port map( A1 => B(11), A2 => n262, ZN => n125);
   U125 : NAND2_X1 port map( A1 => B(10), A2 => n261, ZN => n128);
   U126 : NAND2_X1 port map( A1 => B(18), A2 => n266, ZN => n104);
   U127 : NAND2_X1 port map( A1 => B(14), A2 => n264, ZN => n116);
   U128 : NAND2_X1 port map( A1 => B(5), A2 => n256, ZN => n143);
   U129 : NAND2_X1 port map( A1 => B(7), A2 => n258, ZN => n137);
   U130 : NAND2_X1 port map( A1 => B(27), A2 => n273, ZN => n77);
   U131 : NAND2_X1 port map( A1 => B(23), A2 => n269, ZN => n89);
   U132 : NAND2_X1 port map( A1 => B(25), A2 => n271, ZN => n83);
   U133 : NAND2_X1 port map( A1 => B(15), A2 => n289, ZN => n113);
   U134 : OR2_X1 port map( A1 => n272, A2 => B(26), ZN => n163);
   U135 : OR2_X1 port map( A1 => n257, A2 => B(6), ZN => n193);
   U136 : NAND2_X1 port map( A1 => B(2), A2 => n253, ZN => n153);
   U137 : INV_X1 port map( A => B(31), ZN => n277);
   U138 : AND2_X1 port map( A1 => B(4), A2 => n255, ZN => n147);
   U139 : OR2_X1 port map( A1 => n261, A2 => B(10), ZN => n187);
   U140 : OR2_X1 port map( A1 => n266, A2 => B(18), ZN => n175);
   U141 : OR2_X1 port map( A1 => n264, A2 => B(14), ZN => n181);
   U142 : AND2_X1 port map( A1 => B(12), A2 => n291, ZN => n123);
   U143 : AND2_X1 port map( A1 => B(16), A2 => n288, ZN => n111);
   U144 : INV_X1 port map( A => B(30), ZN => net52651);
   U145 : AND2_X1 port map( A1 => B(20), A2 => n290, ZN => n99);
   U146 : AND2_X1 port map( A1 => B(24), A2 => n270, ZN => n87);
   U147 : INV_X1 port map( A => B(1), ZN => n286);
   U148 : INV_X1 port map( A => n202, ZN => n276);
   U149 : INV_X1 port map( A => A(19), ZN => n287);
   U150 : NOR2_X1 port map( A1 => n277, A2 => A(31), ZN => n66);
   U151 : INV_X1 port map( A => A(16), ZN => n288);
   U152 : INV_X1 port map( A => A(15), ZN => n289);
   U153 : INV_X1 port map( A => A(12), ZN => n291);
   U154 : INV_X1 port map( A => A(20), ZN => n290);
   U155 : NAND2_X1 port map( A1 => A(31), A2 => n277, ZN => n65);
   U156 : INV_X1 port map( A => n150, ZN => n283);
   U157 : OAI211_X1 port map( C1 => A(1), C2 => n212, A => n285, B => n152, ZN 
                           => n199);
   U158 : INV_X1 port map( A => n201, ZN => n285);
   U159 : AOI21_X1 port map( B1 => n200, B2 => A(1), A => n286, ZN => n201);
   U160 : AOI21_X1 port map( B1 => net52652, B2 => n65, A => n66, ZN => n292);
   U161 : NOR2_X1 port map( A1 => n263, A2 => B(13), ZN => n120);
   U162 : AOI21_X1 port map( B1 => n152, B2 => n151, A => n284, ZN => n148);
   U163 : AOI22_X1 port map( A1 => n286, A2 => n154, B1 => n155, B2 => A(1), ZN
                           => n151);
   U164 : AOI21_X1 port map( B1 => n130, B2 => n131, A => n132, ZN => n127);
   U165 : AOI21_X1 port map( B1 => n133, B2 => n134, A => n135, ZN => n130);
   U166 : AOI21_X1 port map( B1 => n136, B2 => n137, A => n138, ZN => n133);
   U167 : OR2_X1 port map( A1 => n268, A2 => B(22), ZN => n169);
   U168 : NAND2_X1 port map( A1 => B(22), A2 => n268, ZN => n92);
   U169 : NOR2_X1 port map( A1 => n274, A2 => B(28), ZN => n162);
   U171 : AND2_X1 port map( A1 => B(28), A2 => n274, ZN => n75);
   U172 : AOI21_X1 port map( B1 => n142, B2 => n143, A => n144, ZN => n139);
   U173 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n145);
   U175 : NAND2_X1 port map( A1 => B(21), A2 => n267, ZN => n95);
   U176 : NOR2_X1 port map( A1 => n267, A2 => B(21), ZN => n96);
   U177 : AND2_X1 port map( A1 => n292, A2 => n276, ZN => EQ);
   U178 : AOI21_X1 port map( B1 => n139, B2 => n281, A => n280, ZN => n136);
   U179 : NOR2_X1 port map( A1 => n252, A2 => B(0), ZN => n200);
   U180 : AOI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n142);
   U181 : NAND2_X1 port map( A1 => B(0), A2 => n252, ZN => n155);
   U182 : NOR2_X1 port map( A1 => n259, A2 => B(8), ZN => n192);
   U183 : AND2_X1 port map( A1 => B(8), A2 => n259, ZN => n135);
   U184 : INV_X1 port map( A => A(0), ZN => n252);
   U185 : INV_X1 port map( A => A(2), ZN => n253);
   U186 : INV_X1 port map( A => A(3), ZN => n254);
   U187 : INV_X1 port map( A => A(4), ZN => n255);
   U188 : INV_X1 port map( A => A(5), ZN => n256);
   U189 : INV_X1 port map( A => A(6), ZN => n257);
   U190 : INV_X1 port map( A => A(7), ZN => n258);
   U191 : INV_X1 port map( A => A(8), ZN => n259);
   U192 : INV_X1 port map( A => A(9), ZN => n260);
   U193 : INV_X1 port map( A => A(10), ZN => n261);
   U194 : INV_X1 port map( A => A(11), ZN => n262);
   U195 : INV_X1 port map( A => A(13), ZN => n263);
   U196 : INV_X1 port map( A => A(14), ZN => n264);
   U197 : INV_X1 port map( A => A(17), ZN => n265);
   U198 : INV_X1 port map( A => A(18), ZN => n266);
   U199 : INV_X1 port map( A => A(21), ZN => n267);
   U200 : INV_X1 port map( A => A(22), ZN => n268);
   U201 : INV_X1 port map( A => A(23), ZN => n269);
   U202 : INV_X1 port map( A => A(24), ZN => n270);
   U203 : INV_X1 port map( A => A(25), ZN => n271);
   U204 : INV_X1 port map( A => A(26), ZN => n272);
   U205 : INV_X1 port map( A => A(27), ZN => n273);
   U206 : INV_X1 port map( A => A(28), ZN => n274);
   U207 : INV_X1 port map( A => A(29), ZN => n275);
   U208 : INV_X1 port map( A => A(30), ZN => net54692);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity SUMGEN_NBIT32_NBLOCKS8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
         std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
         std_logic_vector (31 downto 0));

end SUMGEN_NBIT32_NBLOCKS8_1;

architecture SYN_STRUCTURAL of SUMGEN_NBIT32_NBLOCKS8_1 is

   component CSblock_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082 : std_logic;

begin
   
   block_i_0 : CSblock_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), cin => cin_vect(0), Y(3) => 
                           SUM(3), Y(2) => SUM(2), Y(1) => SUM(1), Y(0) => 
                           SUM(0), Co => n_1076);
   block_i_1 : CSblock_NBIT4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), cin => cin_vect(1), Y(3) => 
                           SUM(7), Y(2) => SUM(6), Y(1) => SUM(5), Y(0) => 
                           SUM(4), Co => n_1077);
   block_i_2 : CSblock_NBIT4_6 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), cin => cin_vect(2), Y(3)
                           => SUM(11), Y(2) => SUM(10), Y(1) => SUM(9), Y(0) =>
                           SUM(8), Co => n_1078);
   block_i_3 : CSblock_NBIT4_5 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), cin => cin_vect(3), 
                           Y(3) => SUM(15), Y(2) => SUM(14), Y(1) => SUM(13), 
                           Y(0) => SUM(12), Co => n_1079);
   block_i_4 : CSblock_NBIT4_4 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), cin => cin_vect(4), 
                           Y(3) => SUM(19), Y(2) => SUM(18), Y(1) => SUM(17), 
                           Y(0) => SUM(16), Co => n_1080);
   block_i_5 : CSblock_NBIT4_3 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), cin => cin_vect(5), 
                           Y(3) => SUM(23), Y(2) => SUM(22), Y(1) => SUM(21), 
                           Y(0) => SUM(20), Co => n_1081);
   block_i_6 : CSblock_NBIT4_2 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), cin => cin_vect(6), 
                           Y(3) => SUM(27), Y(2) => SUM(26), Y(1) => SUM(25), 
                           Y(0) => SUM(24), Co => n_1082);
   block_i_7 : CSblock_NBIT4_1 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), cin => cin_vect(7), 
                           Y(3) => SUM(31), Y(2) => SUM(30), Y(1) => SUM(29), 
                           Y(0) => SUM(28), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   component GENERAL_G_1
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_2
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_3
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_4
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_1
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_2
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_3
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_4
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_5
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_6
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_5
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_7
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_6
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_7
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_8
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_9
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_10
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_11
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_12
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_13
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_14
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_15
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_16
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_17
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_18
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_19
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_20
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_21
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_22
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_23
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_24
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_25
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_26
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_8
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_27
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_9
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_1
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_2
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_3
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_4
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_5
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_6
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_7
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_8
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_9
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_10
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_11
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_12
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_13
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_14
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_15
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_16
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_17
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_18
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_19
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_20
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_21
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_22
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_23
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_24
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_25
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_26
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_27
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_28
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_29
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_30
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_31
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component GENERAL_G_10
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_32
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, first_generate, p_vett_4_3_port, p_vett_4_2_port, 
      p_vett_3_3_port, p_vett_3_2_port, p_vett_3_1_port, p_vett_2_7_port, 
      p_vett_2_6_port, p_vett_2_5_port, p_vett_2_4_port, p_vett_2_3_port, 
      p_vett_2_2_port, p_vett_2_1_port, p_vett_1_15_port, p_vett_1_14_port, 
      p_vett_1_13_port, p_vett_1_12_port, p_vett_1_11_port, p_vett_1_10_port, 
      p_vett_1_9_port, p_vett_1_8_port, p_vett_1_7_port, p_vett_1_6_port, 
      p_vett_1_5_port, p_vett_1_4_port, p_vett_1_3_port, p_vett_1_2_port, 
      p_vett_1_1_port, p_vett_0_31_port, p_vett_0_30_port, p_vett_0_29_port, 
      p_vett_0_28_port, p_vett_0_27_port, p_vett_0_26_port, p_vett_0_25_port, 
      p_vett_0_24_port, p_vett_0_23_port, p_vett_0_22_port, p_vett_0_21_port, 
      p_vett_0_20_port, p_vett_0_19_port, p_vett_0_18_port, p_vett_0_17_port, 
      p_vett_0_16_port, p_vett_0_15_port, p_vett_0_14_port, p_vett_0_13_port, 
      p_vett_0_12_port, p_vett_0_11_port, p_vett_0_10_port, p_vett_0_9_port, 
      p_vett_0_8_port, p_vett_0_7_port, p_vett_0_6_port, p_vett_0_5_port, 
      p_vett_0_4_port, p_vett_0_3_port, p_vett_0_2_port, p_vett_0_1_port, 
      p_vett_0_0_port, g_vett_4_3_port, g_vett_4_2_port, g_vett_3_3_port, 
      g_vett_3_2_port, g_vett_3_1_port, g_vett_2_7_port, g_vett_2_6_port, 
      g_vett_2_5_port, g_vett_2_4_port, g_vett_2_3_port, g_vett_2_2_port, 
      g_vett_2_1_port, g_vett_1_15_port, g_vett_1_14_port, g_vett_1_13_port, 
      g_vett_1_12_port, g_vett_1_11_port, g_vett_1_10_port, g_vett_1_9_port, 
      g_vett_1_8_port, g_vett_1_7_port, g_vett_1_6_port, g_vett_1_5_port, 
      g_vett_1_4_port, g_vett_1_3_port, g_vett_1_2_port, g_vett_1_1_port, 
      g_vett_1_0_port, g_vett_0_31_port, g_vett_0_30_port, g_vett_0_29_port, 
      g_vett_0_28_port, g_vett_0_27_port, g_vett_0_26_port, g_vett_0_25_port, 
      g_vett_0_24_port, g_vett_0_23_port, g_vett_0_22_port, g_vett_0_21_port, 
      g_vett_0_20_port, g_vett_0_19_port, g_vett_0_18_port, g_vett_0_17_port, 
      g_vett_0_16_port, g_vett_0_15_port, g_vett_0_14_port, g_vett_0_13_port, 
      g_vett_0_12_port, g_vett_0_11_port, g_vett_0_10_port, g_vett_0_9_port, 
      g_vett_0_8_port, g_vett_0_7_port, g_vett_0_6_port, g_vett_0_5_port, 
      g_vett_0_4_port, g_vett_0_3_port, g_vett_0_2_port, g_vett_0_1_port, 
      g_vett_0_0_port, n_1083 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Cin );
   
   PGblock_first : PG_block_32 port map( A => A(0), B => B(0), G => 
                           first_generate, P => p_vett_0_0_port);
   G_first : GENERAL_G_10 port map( G_in => first_generate, P_in => 
                           p_vett_0_0_port, G_in_prev => Cin, G_out => 
                           g_vett_0_0_port);
   PG_0_1 : PG_block_31 port map( A => A(1), B => B(1), G => g_vett_0_1_port, P
                           => p_vett_0_1_port);
   PG_0_2 : PG_block_30 port map( A => A(2), B => B(2), G => g_vett_0_2_port, P
                           => p_vett_0_2_port);
   PG_0_3 : PG_block_29 port map( A => A(3), B => B(3), G => g_vett_0_3_port, P
                           => p_vett_0_3_port);
   PG_0_4 : PG_block_28 port map( A => A(4), B => B(4), G => g_vett_0_4_port, P
                           => p_vett_0_4_port);
   PG_0_5 : PG_block_27 port map( A => A(5), B => B(5), G => g_vett_0_5_port, P
                           => p_vett_0_5_port);
   PG_0_6 : PG_block_26 port map( A => A(6), B => B(6), G => g_vett_0_6_port, P
                           => p_vett_0_6_port);
   PG_0_7 : PG_block_25 port map( A => A(7), B => B(7), G => g_vett_0_7_port, P
                           => p_vett_0_7_port);
   PG_0_8 : PG_block_24 port map( A => A(8), B => B(8), G => g_vett_0_8_port, P
                           => p_vett_0_8_port);
   PG_0_9 : PG_block_23 port map( A => A(9), B => B(9), G => g_vett_0_9_port, P
                           => p_vett_0_9_port);
   PG_0_10 : PG_block_22 port map( A => A(10), B => B(10), G => 
                           g_vett_0_10_port, P => p_vett_0_10_port);
   PG_0_11 : PG_block_21 port map( A => A(11), B => B(11), G => 
                           g_vett_0_11_port, P => p_vett_0_11_port);
   PG_0_12 : PG_block_20 port map( A => A(12), B => B(12), G => 
                           g_vett_0_12_port, P => p_vett_0_12_port);
   PG_0_13 : PG_block_19 port map( A => A(13), B => B(13), G => 
                           g_vett_0_13_port, P => p_vett_0_13_port);
   PG_0_14 : PG_block_18 port map( A => A(14), B => B(14), G => 
                           g_vett_0_14_port, P => p_vett_0_14_port);
   PG_0_15 : PG_block_17 port map( A => A(15), B => B(15), G => 
                           g_vett_0_15_port, P => p_vett_0_15_port);
   PG_0_16 : PG_block_16 port map( A => A(16), B => B(16), G => 
                           g_vett_0_16_port, P => p_vett_0_16_port);
   PG_0_17 : PG_block_15 port map( A => A(17), B => B(17), G => 
                           g_vett_0_17_port, P => p_vett_0_17_port);
   PG_0_18 : PG_block_14 port map( A => A(18), B => B(18), G => 
                           g_vett_0_18_port, P => p_vett_0_18_port);
   PG_0_19 : PG_block_13 port map( A => A(19), B => B(19), G => 
                           g_vett_0_19_port, P => p_vett_0_19_port);
   PG_0_20 : PG_block_12 port map( A => A(20), B => B(20), G => 
                           g_vett_0_20_port, P => p_vett_0_20_port);
   PG_0_21 : PG_block_11 port map( A => A(21), B => B(21), G => 
                           g_vett_0_21_port, P => p_vett_0_21_port);
   PG_0_22 : PG_block_10 port map( A => A(22), B => B(22), G => 
                           g_vett_0_22_port, P => p_vett_0_22_port);
   PG_0_23 : PG_block_9 port map( A => A(23), B => B(23), G => g_vett_0_23_port
                           , P => p_vett_0_23_port);
   PG_0_24 : PG_block_8 port map( A => A(24), B => B(24), G => g_vett_0_24_port
                           , P => p_vett_0_24_port);
   PG_0_25 : PG_block_7 port map( A => A(25), B => B(25), G => g_vett_0_25_port
                           , P => p_vett_0_25_port);
   PG_0_26 : PG_block_6 port map( A => A(26), B => B(26), G => g_vett_0_26_port
                           , P => p_vett_0_26_port);
   PG_0_27 : PG_block_5 port map( A => A(27), B => B(27), G => g_vett_0_27_port
                           , P => p_vett_0_27_port);
   PG_0_28 : PG_block_4 port map( A => A(28), B => B(28), G => g_vett_0_28_port
                           , P => p_vett_0_28_port);
   PG_0_29 : PG_block_3 port map( A => A(29), B => B(29), G => g_vett_0_29_port
                           , P => p_vett_0_29_port);
   PG_0_30 : PG_block_2 port map( A => A(30), B => B(30), G => g_vett_0_30_port
                           , P => p_vett_0_30_port);
   PG_0_31 : PG_block_1 port map( A => A(31), B => B(31), G => g_vett_0_31_port
                           , P => p_vett_0_31_port);
   G_0_0_0 : GENERAL_G_9 port map( G_in => g_vett_0_1_port, P_in => 
                           p_vett_0_1_port, G_in_prev => g_vett_0_0_port, G_out
                           => g_vett_1_0_port);
   PG_1_0_0 : GENERAL_PG_27 port map( G_in => g_vett_0_3_port, P_in => 
                           p_vett_0_3_port, G_in_prev => g_vett_0_2_port, 
                           P_in_prev => p_vett_0_2_port, G_out => 
                           g_vett_1_1_port, P_out => p_vett_1_1_port);
   G_1_0_0 : GENERAL_G_8 port map( G_in => g_vett_1_1_port, P_in => 
                           p_vett_1_1_port, G_in_prev => g_vett_1_0_port, G_out
                           => Co_1_port);
   PG_2_0_1 : GENERAL_PG_26 port map( G_in => g_vett_0_5_port, P_in => 
                           p_vett_0_5_port, G_in_prev => g_vett_0_4_port, 
                           P_in_prev => p_vett_0_4_port, G_out => 
                           g_vett_1_2_port, P_out => p_vett_1_2_port);
   PG_3_0_1 : GENERAL_PG_25 port map( G_in => g_vett_0_7_port, P_in => 
                           p_vett_0_7_port, G_in_prev => g_vett_0_6_port, 
                           P_in_prev => p_vett_0_6_port, G_out => 
                           g_vett_1_3_port, P_out => p_vett_1_3_port);
   PG_4_0_1 : GENERAL_PG_24 port map( G_in => g_vett_1_3_port, P_in => 
                           p_vett_1_3_port, G_in_prev => g_vett_1_2_port, 
                           P_in_prev => p_vett_1_2_port, G_out => 
                           g_vett_2_1_port, P_out => p_vett_2_1_port);
   PG_2_0_2 : GENERAL_PG_23 port map( G_in => g_vett_0_9_port, P_in => 
                           p_vett_0_9_port, G_in_prev => g_vett_0_8_port, 
                           P_in_prev => p_vett_0_8_port, G_out => 
                           g_vett_1_4_port, P_out => p_vett_1_4_port);
   PG_3_0_2 : GENERAL_PG_22 port map( G_in => g_vett_0_11_port, P_in => 
                           p_vett_0_11_port, G_in_prev => g_vett_0_10_port, 
                           P_in_prev => p_vett_0_10_port, G_out => 
                           g_vett_1_5_port, P_out => p_vett_1_5_port);
   PG_4_0_2 : GENERAL_PG_21 port map( G_in => g_vett_1_5_port, P_in => 
                           p_vett_1_5_port, G_in_prev => g_vett_1_4_port, 
                           P_in_prev => p_vett_1_4_port, G_out => 
                           g_vett_2_2_port, P_out => p_vett_2_2_port);
   PG_2_0_3 : GENERAL_PG_20 port map( G_in => g_vett_0_13_port, P_in => 
                           p_vett_0_13_port, G_in_prev => g_vett_0_12_port, 
                           P_in_prev => p_vett_0_12_port, G_out => 
                           g_vett_1_6_port, P_out => p_vett_1_6_port);
   PG_3_0_3 : GENERAL_PG_19 port map( G_in => g_vett_0_15_port, P_in => 
                           p_vett_0_15_port, G_in_prev => g_vett_0_14_port, 
                           P_in_prev => p_vett_0_14_port, G_out => 
                           g_vett_1_7_port, P_out => p_vett_1_7_port);
   PG_4_0_3 : GENERAL_PG_18 port map( G_in => g_vett_1_7_port, P_in => 
                           p_vett_1_7_port, G_in_prev => g_vett_1_6_port, 
                           P_in_prev => p_vett_1_6_port, G_out => 
                           g_vett_2_3_port, P_out => p_vett_2_3_port);
   PG_2_0_4 : GENERAL_PG_17 port map( G_in => g_vett_0_17_port, P_in => 
                           p_vett_0_17_port, G_in_prev => g_vett_0_16_port, 
                           P_in_prev => p_vett_0_16_port, G_out => 
                           g_vett_1_8_port, P_out => p_vett_1_8_port);
   PG_3_0_4 : GENERAL_PG_16 port map( G_in => g_vett_0_19_port, P_in => 
                           p_vett_0_19_port, G_in_prev => g_vett_0_18_port, 
                           P_in_prev => p_vett_0_18_port, G_out => 
                           g_vett_1_9_port, P_out => p_vett_1_9_port);
   PG_4_0_4 : GENERAL_PG_15 port map( G_in => g_vett_1_9_port, P_in => 
                           p_vett_1_9_port, G_in_prev => g_vett_1_8_port, 
                           P_in_prev => p_vett_1_8_port, G_out => 
                           g_vett_2_4_port, P_out => p_vett_2_4_port);
   PG_2_0_5 : GENERAL_PG_14 port map( G_in => g_vett_0_21_port, P_in => 
                           p_vett_0_21_port, G_in_prev => g_vett_0_20_port, 
                           P_in_prev => p_vett_0_20_port, G_out => 
                           g_vett_1_10_port, P_out => p_vett_1_10_port);
   PG_3_0_5 : GENERAL_PG_13 port map( G_in => g_vett_0_23_port, P_in => 
                           p_vett_0_23_port, G_in_prev => g_vett_0_22_port, 
                           P_in_prev => p_vett_0_22_port, G_out => 
                           g_vett_1_11_port, P_out => p_vett_1_11_port);
   PG_4_0_5 : GENERAL_PG_12 port map( G_in => g_vett_1_11_port, P_in => 
                           p_vett_1_11_port, G_in_prev => g_vett_1_10_port, 
                           P_in_prev => p_vett_1_10_port, G_out => 
                           g_vett_2_5_port, P_out => p_vett_2_5_port);
   PG_2_0_6 : GENERAL_PG_11 port map( G_in => g_vett_0_25_port, P_in => 
                           p_vett_0_25_port, G_in_prev => g_vett_0_24_port, 
                           P_in_prev => p_vett_0_24_port, G_out => 
                           g_vett_1_12_port, P_out => p_vett_1_12_port);
   PG_3_0_6 : GENERAL_PG_10 port map( G_in => g_vett_0_27_port, P_in => 
                           p_vett_0_27_port, G_in_prev => g_vett_0_26_port, 
                           P_in_prev => p_vett_0_26_port, G_out => 
                           g_vett_1_13_port, P_out => p_vett_1_13_port);
   PG_4_0_6 : GENERAL_PG_9 port map( G_in => g_vett_1_13_port, P_in => 
                           p_vett_1_13_port, G_in_prev => g_vett_1_12_port, 
                           P_in_prev => p_vett_1_12_port, G_out => 
                           g_vett_2_6_port, P_out => p_vett_2_6_port);
   PG_2_0_7 : GENERAL_PG_8 port map( G_in => g_vett_0_29_port, P_in => 
                           p_vett_0_29_port, G_in_prev => g_vett_0_28_port, 
                           P_in_prev => p_vett_0_28_port, G_out => 
                           g_vett_1_14_port, P_out => p_vett_1_14_port);
   PG_3_0_7 : GENERAL_PG_7 port map( G_in => g_vett_0_31_port, P_in => 
                           p_vett_0_31_port, G_in_prev => g_vett_0_30_port, 
                           P_in_prev => p_vett_0_30_port, G_out => 
                           g_vett_1_15_port, P_out => p_vett_1_15_port);
   PG_4_0_7 : GENERAL_PG_6 port map( G_in => g_vett_1_15_port, P_in => 
                           p_vett_1_15_port, G_in_prev => g_vett_1_14_port, 
                           P_in_prev => p_vett_1_14_port, G_out => 
                           g_vett_2_7_port, P_out => p_vett_2_7_port);
   G_2_1_0 : GENERAL_G_7 port map( G_in => g_vett_2_1_port, P_in => 
                           p_vett_2_1_port, G_in_prev => Co_1_port, G_out => 
                           Co_2_port);
   PG_5_1_0 : GENERAL_PG_5 port map( G_in => g_vett_2_3_port, P_in => 
                           p_vett_2_3_port, G_in_prev => g_vett_2_2_port, 
                           P_in_prev => p_vett_2_2_port, G_out => 
                           g_vett_3_1_port, P_out => p_vett_3_1_port);
   G_3_1_0 : GENERAL_G_6 port map( G_in => g_vett_2_2_port, P_in => 
                           p_vett_2_2_port, G_in_prev => Co_2_port, G_out => 
                           Co_3_port);
   G_4_1_0 : GENERAL_G_5 port map( G_in => g_vett_3_1_port, P_in => 
                           p_vett_3_1_port, G_in_prev => Co_2_port, G_out => 
                           Co_4_port);
   PG_6_1_1 : GENERAL_PG_4 port map( G_in => g_vett_2_5_port, P_in => 
                           p_vett_2_5_port, G_in_prev => g_vett_2_4_port, 
                           P_in_prev => p_vett_2_4_port, G_out => 
                           g_vett_3_2_port, P_out => p_vett_3_2_port);
   PG_7_1_1 : GENERAL_PG_3 port map( G_in => g_vett_2_7_port, P_in => 
                           p_vett_2_7_port, G_in_prev => g_vett_2_6_port, 
                           P_in_prev => p_vett_2_6_port, G_out => 
                           g_vett_3_3_port, P_out => p_vett_3_3_port);
   PG_8_1_1 : GENERAL_PG_2 port map( G_in => g_vett_2_6_port, P_in => 
                           p_vett_2_6_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_2_port, P_out => p_vett_4_2_port);
   PG_9_1_1 : GENERAL_PG_1 port map( G_in => g_vett_3_3_port, P_in => 
                           p_vett_3_3_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_3_port, P_out => p_vett_4_3_port);
   G_5_2_0 : GENERAL_G_4 port map( G_in => g_vett_2_4_port, P_in => 
                           p_vett_2_4_port, G_in_prev => Co_4_port, G_out => 
                           Co_5_port);
   G_6_2_1 : GENERAL_G_3 port map( G_in => g_vett_3_2_port, P_in => 
                           p_vett_3_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_6_port);
   G_7_2_2 : GENERAL_G_2 port map( G_in => g_vett_4_2_port, P_in => 
                           p_vett_4_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_7_port);
   G_8_2_3 : GENERAL_G_1 port map( G_in => g_vett_4_3_port, P_in => 
                           p_vett_4_3_port, G_in_prev => Co_4_port, G_out => 
                           n_1083);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_25;

architecture SYN_structural of CSblock_NBIT4_25 is

   component MUX21_GENERIC_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1084, n_1085, n_1086 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_50 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_49 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_50 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_49 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1084, Y(2) => 
                           n_1085, Y(1) => n_1086, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_26;

architecture SYN_structural of CSblock_NBIT4_26 is

   component MUX21_GENERIC_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1087, n_1088, n_1089 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_52 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_51 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_52 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_51 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1087, Y(2) => 
                           n_1088, Y(1) => n_1089, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_27;

architecture SYN_structural of CSblock_NBIT4_27 is

   component MUX21_GENERIC_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1090, n_1091, n_1092 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_54 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_53 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_54 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_53 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1090, Y(2) => 
                           n_1091, Y(1) => n_1092, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_28;

architecture SYN_structural of CSblock_NBIT4_28 is

   component MUX21_GENERIC_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1093, n_1094, n_1095 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_55 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_56 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_55 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1093, Y(2) => 
                           n_1094, Y(1) => n_1095, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_29;

architecture SYN_structural of CSblock_NBIT4_29 is

   component MUX21_GENERIC_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1096, n_1097, n_1098 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_58 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_57 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_58 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_57 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1096, Y(2) => 
                           n_1097, Y(1) => n_1098, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_30;

architecture SYN_structural of CSblock_NBIT4_30 is

   component MUX21_GENERIC_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1099, n_1100, n_1101 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_60 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_59 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_60 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_59 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1099, Y(2) => 
                           n_1100, Y(1) => n_1101, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_31;

architecture SYN_structural of CSblock_NBIT4_31 is

   component MUX21_GENERIC_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1102, n_1103, n_1104 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_62 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_61 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_62 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_61 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1102, Y(2) => 
                           n_1103, Y(1) => n_1104, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CSblock_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  Co : out std_logic);

end CSblock_NBIT4_0;

architecture SYN_structural of CSblock_NBIT4_0 is

   component MUX21_GENERIC_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, out0_0_port, 
      cout0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, 
      cout1_0_port, n_1105, n_1106, n_1107 : std_logic;

begin
   
   X_Logic0_port <= '0';
   add0 : RCA_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out0_3_port, S(2) => out0_2_port, S(1) => 
                           out0_1_port, S(0) => out0_0_port, Co => cout0_0_port
                           );
   add1 : RCA_NBIT4_63 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out1_3_port, S(2) => out1_2_port, S(1) => 
                           out1_1_port, S(0) => out1_0_port, Co => cout1_0_port
                           );
   muxSum : MUX21_GENERIC_NBIT4_0 port map( A(3) => out0_3_port, A(2) => 
                           out0_2_port, A(1) => out0_1_port, A(0) => 
                           out0_0_port, B(3) => out1_3_port, B(2) => 
                           out1_2_port, B(1) => out1_1_port, B(0) => 
                           out1_0_port, SEL => cin, Y(3) => Y(3), Y(2) => Y(2),
                           Y(1) => Y(1), Y(0) => Y(0));
   muxCout : MUX21_GENERIC_NBIT4_63 port map( A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           cout0_0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           cout1_0_port, SEL => cin, Y(3) => n_1105, Y(2) => 
                           n_1106, Y(1) => n_1107, Y(0) => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_31 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_31;

architecture SYN_BEHAVIORAL of GENERAL_G_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_32 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_32;

architecture SYN_BEHAVIORAL of GENERAL_G_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_33 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_33;

architecture SYN_BEHAVIORAL of GENERAL_G_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_34 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_34;

architecture SYN_BEHAVIORAL of GENERAL_G_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_82 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_82;

architecture SYN_BEHAVIORAL of GENERAL_PG_82 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_83 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_83;

architecture SYN_BEHAVIORAL of GENERAL_PG_83 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_84 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_84;

architecture SYN_BEHAVIORAL of GENERAL_PG_84 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_85 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_85;

architecture SYN_BEHAVIORAL of GENERAL_PG_85 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_35 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_35;

architecture SYN_BEHAVIORAL of GENERAL_G_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_36 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_36;

architecture SYN_BEHAVIORAL of GENERAL_G_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_86 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_86;

architecture SYN_BEHAVIORAL of GENERAL_PG_86 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_37 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_37;

architecture SYN_BEHAVIORAL of GENERAL_G_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_87 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_87;

architecture SYN_BEHAVIORAL of GENERAL_PG_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_88 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_88;

architecture SYN_BEHAVIORAL of GENERAL_PG_88 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_89 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_89;

architecture SYN_BEHAVIORAL of GENERAL_PG_89 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_90 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_90;

architecture SYN_BEHAVIORAL of GENERAL_PG_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_91 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_91;

architecture SYN_BEHAVIORAL of GENERAL_PG_91 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_92 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_92;

architecture SYN_BEHAVIORAL of GENERAL_PG_92 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_93 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_93;

architecture SYN_BEHAVIORAL of GENERAL_PG_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_94 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_94;

architecture SYN_BEHAVIORAL of GENERAL_PG_94 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_95 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_95;

architecture SYN_BEHAVIORAL of GENERAL_PG_95 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_96 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_96;

architecture SYN_BEHAVIORAL of GENERAL_PG_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_97 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_97;

architecture SYN_BEHAVIORAL of GENERAL_PG_97 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_98 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_98;

architecture SYN_BEHAVIORAL of GENERAL_PG_98 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_99 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_99;

architecture SYN_BEHAVIORAL of GENERAL_PG_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_100 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_100;

architecture SYN_BEHAVIORAL of GENERAL_PG_100 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_101 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_101;

architecture SYN_BEHAVIORAL of GENERAL_PG_101 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n4, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_102 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_102;

architecture SYN_BEHAVIORAL of GENERAL_PG_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_103 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_103;

architecture SYN_BEHAVIORAL of GENERAL_PG_103 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_104 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_104;

architecture SYN_BEHAVIORAL of GENERAL_PG_104 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_105 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_105;

architecture SYN_BEHAVIORAL of GENERAL_PG_105 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_106 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_106;

architecture SYN_BEHAVIORAL of GENERAL_PG_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);
   U3 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_107 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_107;

architecture SYN_BEHAVIORAL of GENERAL_PG_107 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_38 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_38;

architecture SYN_BEHAVIORAL of GENERAL_G_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_PG_0 is

   port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : out 
         std_logic);

end GENERAL_PG_0;

architecture SYN_BEHAVIORAL of GENERAL_PG_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_in_prev, A2 => P_in, ZN => P_out);
   U2 : INV_X1 port map( A => n2, ZN => G_out);
   U3 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_39 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_39;

architecture SYN_BEHAVIORAL of GENERAL_G_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => G_out);
   U2 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_97 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_97;

architecture SYN_BEHAVIORAL of PG_block_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_98 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_98;

architecture SYN_BEHAVIORAL of PG_block_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_99 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_99;

architecture SYN_BEHAVIORAL of PG_block_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_100 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_100;

architecture SYN_BEHAVIORAL of PG_block_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_101 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_101;

architecture SYN_BEHAVIORAL of PG_block_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_102 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_102;

architecture SYN_BEHAVIORAL of PG_block_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_103 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_103;

architecture SYN_BEHAVIORAL of PG_block_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_104 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_104;

architecture SYN_BEHAVIORAL of PG_block_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_105 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_105;

architecture SYN_BEHAVIORAL of PG_block_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_106 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_106;

architecture SYN_BEHAVIORAL of PG_block_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_107 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_107;

architecture SYN_BEHAVIORAL of PG_block_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_108 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_108;

architecture SYN_BEHAVIORAL of PG_block_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_109 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_109;

architecture SYN_BEHAVIORAL of PG_block_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_110 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_110;

architecture SYN_BEHAVIORAL of PG_block_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_111 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_111;

architecture SYN_BEHAVIORAL of PG_block_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_112 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_112;

architecture SYN_BEHAVIORAL of PG_block_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_113 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_113;

architecture SYN_BEHAVIORAL of PG_block_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_114 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_114;

architecture SYN_BEHAVIORAL of PG_block_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_115 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_115;

architecture SYN_BEHAVIORAL of PG_block_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_116 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_116;

architecture SYN_BEHAVIORAL of PG_block_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_117 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_117;

architecture SYN_BEHAVIORAL of PG_block_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_118 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_118;

architecture SYN_BEHAVIORAL of PG_block_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_119 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_119;

architecture SYN_BEHAVIORAL of PG_block_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_120 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_120;

architecture SYN_BEHAVIORAL of PG_block_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_121 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_121;

architecture SYN_BEHAVIORAL of PG_block_121 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_122 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_122;

architecture SYN_BEHAVIORAL of PG_block_122 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_123 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_123;

architecture SYN_BEHAVIORAL of PG_block_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_124 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_124;

architecture SYN_BEHAVIORAL of PG_block_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_125 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_125;

architecture SYN_BEHAVIORAL of PG_block_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_126 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_126;

architecture SYN_BEHAVIORAL of PG_block_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_127 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_127;

architecture SYN_BEHAVIORAL of PG_block_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity GENERAL_G_0 is

   port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);

end GENERAL_G_0;

architecture SYN_BEHAVIORAL of GENERAL_G_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => P_in, B2 => G_in_prev, A => G_in, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => G_out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity PG_block_0 is

   port( A, B : in std_logic;  G, P : out std_logic);

end PG_block_0;

architecture SYN_BEHAVIORAL of PG_block_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n78, ZN => n68);
   U2 : INV_X1 port map( A => n78, ZN => n69);
   U3 : BUF_X1 port map( A => n33, Z => n70);
   U4 : BUF_X1 port map( A => n67, Z => n76);
   U5 : BUF_X1 port map( A => n66, Z => n75);
   U6 : BUF_X1 port map( A => n66, Z => n73);
   U7 : BUF_X1 port map( A => n33, Z => n72);
   U8 : BUF_X1 port map( A => n66, Z => n74);
   U9 : BUF_X1 port map( A => n33, Z => n71);
   U10 : BUF_X1 port map( A => n67, Z => n78);
   U11 : BUF_X1 port map( A => n67, Z => n77);
   U12 : BUF_X1 port map( A => SEL, Z => n67);
   U13 : BUF_X1 port map( A => SEL, Z => n66);
   U14 : BUF_X1 port map( A => SEL, Z => n33);
   U15 : INV_X1 port map( A => n142, ZN => Y(9));
   U16 : AOI22_X1 port map( A1 => A(9), A2 => n68, B1 => n77, B2 => B(9), ZN =>
                           n142);
   U17 : INV_X1 port map( A => n111, ZN => Y(0));
   U18 : AOI22_X1 port map( A1 => A(0), A2 => n68, B1 => B(0), B2 => n77, ZN =>
                           n111);
   U19 : INV_X1 port map( A => n122, ZN => Y(1));
   U20 : AOI22_X1 port map( A1 => A(1), A2 => n68, B1 => B(1), B2 => n74, ZN =>
                           n122);
   U21 : INV_X1 port map( A => n133, ZN => Y(2));
   U22 : AOI22_X1 port map( A1 => A(2), A2 => n69, B1 => B(2), B2 => n71, ZN =>
                           n133);
   U23 : INV_X1 port map( A => n136, ZN => Y(3));
   U24 : AOI22_X1 port map( A1 => A(3), A2 => n69, B1 => B(3), B2 => n71, ZN =>
                           n136);
   U25 : INV_X1 port map( A => n137, ZN => Y(4));
   U26 : AOI22_X1 port map( A1 => A(4), A2 => n68, B1 => B(4), B2 => n71, ZN =>
                           n137);
   U27 : INV_X1 port map( A => n138, ZN => Y(5));
   U28 : AOI22_X1 port map( A1 => A(5), A2 => n69, B1 => B(5), B2 => n70, ZN =>
                           n138);
   U29 : INV_X1 port map( A => n139, ZN => Y(6));
   U30 : AOI22_X1 port map( A1 => A(6), A2 => n68, B1 => B(6), B2 => n70, ZN =>
                           n139);
   U31 : INV_X1 port map( A => n140, ZN => Y(7));
   U32 : AOI22_X1 port map( A1 => A(7), A2 => n69, B1 => B(7), B2 => n70, ZN =>
                           n140);
   U33 : INV_X1 port map( A => n141, ZN => Y(8));
   U34 : AOI22_X1 port map( A1 => A(8), A2 => n68, B1 => B(8), B2 => n70, ZN =>
                           n141);
   U35 : INV_X1 port map( A => n112, ZN => Y(10));
   U36 : AOI22_X1 port map( A1 => A(10), A2 => n68, B1 => B(10), B2 => n77, ZN 
                           => n112);
   U37 : INV_X1 port map( A => n113, ZN => Y(11));
   U38 : AOI22_X1 port map( A1 => A(11), A2 => n68, B1 => B(11), B2 => n77, ZN 
                           => n113);
   U39 : INV_X1 port map( A => n114, ZN => Y(12));
   U40 : AOI22_X1 port map( A1 => A(12), A2 => n68, B1 => B(12), B2 => n76, ZN 
                           => n114);
   U41 : INV_X1 port map( A => n115, ZN => Y(13));
   U42 : AOI22_X1 port map( A1 => A(13), A2 => n68, B1 => B(13), B2 => n76, ZN 
                           => n115);
   U43 : INV_X1 port map( A => n116, ZN => Y(14));
   U44 : AOI22_X1 port map( A1 => A(14), A2 => n68, B1 => B(14), B2 => n76, ZN 
                           => n116);
   U45 : INV_X1 port map( A => n117, ZN => Y(15));
   U46 : AOI22_X1 port map( A1 => A(15), A2 => n68, B1 => B(15), B2 => n76, ZN 
                           => n117);
   U47 : INV_X1 port map( A => n118, ZN => Y(16));
   U48 : AOI22_X1 port map( A1 => A(16), A2 => n68, B1 => B(16), B2 => n75, ZN 
                           => n118);
   U49 : INV_X1 port map( A => n119, ZN => Y(17));
   U50 : AOI22_X1 port map( A1 => A(17), A2 => n68, B1 => B(17), B2 => n75, ZN 
                           => n119);
   U51 : INV_X1 port map( A => n120, ZN => Y(18));
   U52 : AOI22_X1 port map( A1 => A(18), A2 => n68, B1 => B(18), B2 => n75, ZN 
                           => n120);
   U53 : INV_X1 port map( A => n121, ZN => Y(19));
   U54 : AOI22_X1 port map( A1 => A(19), A2 => n68, B1 => B(19), B2 => n75, ZN 
                           => n121);
   U55 : INV_X1 port map( A => n123, ZN => Y(20));
   U56 : AOI22_X1 port map( A1 => A(20), A2 => n69, B1 => B(20), B2 => n74, ZN 
                           => n123);
   U57 : INV_X1 port map( A => n124, ZN => Y(21));
   U58 : AOI22_X1 port map( A1 => A(21), A2 => n69, B1 => B(21), B2 => n74, ZN 
                           => n124);
   U59 : INV_X1 port map( A => n125, ZN => Y(22));
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n69, B1 => B(22), B2 => n73, ZN 
                           => n125);
   U61 : INV_X1 port map( A => n126, ZN => Y(23));
   U62 : AOI22_X1 port map( A1 => A(23), A2 => n69, B1 => B(23), B2 => n73, ZN 
                           => n126);
   U63 : INV_X1 port map( A => n127, ZN => Y(24));
   U64 : AOI22_X1 port map( A1 => A(24), A2 => n69, B1 => B(24), B2 => n73, ZN 
                           => n127);
   U65 : INV_X1 port map( A => n128, ZN => Y(25));
   U66 : AOI22_X1 port map( A1 => A(25), A2 => n69, B1 => B(25), B2 => n73, ZN 
                           => n128);
   U67 : INV_X1 port map( A => n129, ZN => Y(26));
   U68 : AOI22_X1 port map( A1 => A(26), A2 => n69, B1 => B(26), B2 => n72, ZN 
                           => n129);
   U69 : INV_X1 port map( A => n130, ZN => Y(27));
   U70 : AOI22_X1 port map( A1 => A(27), A2 => n69, B1 => B(27), B2 => n72, ZN 
                           => n130);
   U71 : INV_X1 port map( A => n131, ZN => Y(28));
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n69, B1 => B(28), B2 => n72, ZN 
                           => n131);
   U73 : INV_X1 port map( A => n132, ZN => Y(29));
   U74 : AOI22_X1 port map( A1 => A(29), A2 => n69, B1 => B(29), B2 => n72, ZN 
                           => n132);
   U75 : INV_X1 port map( A => n134, ZN => Y(30));
   U76 : AOI22_X1 port map( A1 => A(30), A2 => n69, B1 => B(30), B2 => n74, ZN 
                           => n134);
   U77 : INV_X1 port map( A => n135, ZN => Y(31));
   U78 : AOI22_X1 port map( A1 => A(31), A2 => n69, B1 => B(31), B2 => n71, ZN 
                           => n135);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity SUMGEN_NBIT32_NBLOCKS8_2 is

   port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
         std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
         std_logic_vector (31 downto 0));

end SUMGEN_NBIT32_NBLOCKS8_2;

architecture SYN_STRUCTURAL of SUMGEN_NBIT32_NBLOCKS8_2 is

   component CSblock_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114 : std_logic;

begin
   
   block_i_0 : CSblock_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), cin => cin_vect(0), Y(3) => 
                           SUM(3), Y(2) => SUM(2), Y(1) => SUM(1), Y(0) => 
                           SUM(0), Co => n_1108);
   block_i_1 : CSblock_NBIT4_15 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), cin => cin_vect(1), Y(3) => 
                           SUM(7), Y(2) => SUM(6), Y(1) => SUM(5), Y(0) => 
                           SUM(4), Co => n_1109);
   block_i_2 : CSblock_NBIT4_14 port map( A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), cin => cin_vect(2), Y(3)
                           => SUM(11), Y(2) => SUM(10), Y(1) => SUM(9), Y(0) =>
                           SUM(8), Co => n_1110);
   block_i_3 : CSblock_NBIT4_13 port map( A(3) => A(15), A(2) => A(14), A(1) =>
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), cin => cin_vect(3), 
                           Y(3) => SUM(15), Y(2) => SUM(14), Y(1) => SUM(13), 
                           Y(0) => SUM(12), Co => n_1111);
   block_i_4 : CSblock_NBIT4_12 port map( A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), cin => cin_vect(4), 
                           Y(3) => SUM(19), Y(2) => SUM(18), Y(1) => SUM(17), 
                           Y(0) => SUM(16), Co => n_1112);
   block_i_5 : CSblock_NBIT4_11 port map( A(3) => A(23), A(2) => A(22), A(1) =>
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), cin => cin_vect(5), 
                           Y(3) => SUM(23), Y(2) => SUM(22), Y(1) => SUM(21), 
                           Y(0) => SUM(20), Co => n_1113);
   block_i_6 : CSblock_NBIT4_10 port map( A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), cin => cin_vect(6), 
                           Y(3) => SUM(27), Y(2) => SUM(26), Y(1) => SUM(25), 
                           Y(0) => SUM(24), Co => n_1114);
   block_i_7 : CSblock_NBIT4_9 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), cin => cin_vect(7), 
                           Y(3) => SUM(31), Y(2) => SUM(30), Y(1) => SUM(29), 
                           Y(0) => SUM(28), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 is

   component GENERAL_G_11
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_12
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_13
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_14
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_28
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_29
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_30
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_31
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_15
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_16
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_32
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_17
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_33
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_34
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_35
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_36
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_37
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_38
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_39
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_40
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_41
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_42
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_43
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_44
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_45
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_46
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_47
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_48
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_49
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_50
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_51
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_52
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_53
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_18
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_54
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_19
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_33
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_34
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_35
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_36
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_37
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_38
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_39
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_40
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_41
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_42
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_43
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_44
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_45
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_46
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_47
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_48
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_49
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_50
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_51
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_52
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_53
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_54
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_55
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_56
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_57
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_58
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_59
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_60
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_61
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_62
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_63
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component GENERAL_G_20
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_64
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, first_generate, p_vett_4_3_port, p_vett_4_2_port, 
      p_vett_3_3_port, p_vett_3_2_port, p_vett_3_1_port, p_vett_2_7_port, 
      p_vett_2_6_port, p_vett_2_5_port, p_vett_2_4_port, p_vett_2_3_port, 
      p_vett_2_2_port, p_vett_2_1_port, p_vett_1_15_port, p_vett_1_14_port, 
      p_vett_1_13_port, p_vett_1_12_port, p_vett_1_11_port, p_vett_1_10_port, 
      p_vett_1_9_port, p_vett_1_8_port, p_vett_1_7_port, p_vett_1_6_port, 
      p_vett_1_5_port, p_vett_1_4_port, p_vett_1_3_port, p_vett_1_2_port, 
      p_vett_1_1_port, p_vett_0_31_port, p_vett_0_30_port, p_vett_0_29_port, 
      p_vett_0_28_port, p_vett_0_27_port, p_vett_0_26_port, p_vett_0_25_port, 
      p_vett_0_24_port, p_vett_0_23_port, p_vett_0_22_port, p_vett_0_21_port, 
      p_vett_0_20_port, p_vett_0_19_port, p_vett_0_18_port, p_vett_0_17_port, 
      p_vett_0_16_port, p_vett_0_15_port, p_vett_0_14_port, p_vett_0_13_port, 
      p_vett_0_12_port, p_vett_0_11_port, p_vett_0_10_port, p_vett_0_9_port, 
      p_vett_0_8_port, p_vett_0_7_port, p_vett_0_6_port, p_vett_0_5_port, 
      p_vett_0_4_port, p_vett_0_3_port, p_vett_0_2_port, p_vett_0_1_port, 
      p_vett_0_0_port, g_vett_4_3_port, g_vett_4_2_port, g_vett_3_3_port, 
      g_vett_3_2_port, g_vett_3_1_port, g_vett_2_7_port, g_vett_2_6_port, 
      g_vett_2_5_port, g_vett_2_4_port, g_vett_2_3_port, g_vett_2_2_port, 
      g_vett_2_1_port, g_vett_1_15_port, g_vett_1_14_port, g_vett_1_13_port, 
      g_vett_1_12_port, g_vett_1_11_port, g_vett_1_10_port, g_vett_1_9_port, 
      g_vett_1_8_port, g_vett_1_7_port, g_vett_1_6_port, g_vett_1_5_port, 
      g_vett_1_4_port, g_vett_1_3_port, g_vett_1_2_port, g_vett_1_1_port, 
      g_vett_1_0_port, g_vett_0_31_port, g_vett_0_30_port, g_vett_0_29_port, 
      g_vett_0_28_port, g_vett_0_27_port, g_vett_0_26_port, g_vett_0_25_port, 
      g_vett_0_24_port, g_vett_0_23_port, g_vett_0_22_port, g_vett_0_21_port, 
      g_vett_0_20_port, g_vett_0_19_port, g_vett_0_18_port, g_vett_0_17_port, 
      g_vett_0_16_port, g_vett_0_15_port, g_vett_0_14_port, g_vett_0_13_port, 
      g_vett_0_12_port, g_vett_0_11_port, g_vett_0_10_port, g_vett_0_9_port, 
      g_vett_0_8_port, g_vett_0_7_port, g_vett_0_6_port, g_vett_0_5_port, 
      g_vett_0_4_port, g_vett_0_3_port, g_vett_0_2_port, g_vett_0_1_port, 
      g_vett_0_0_port, n_1115 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Cin );
   
   PGblock_first : PG_block_64 port map( A => A(0), B => B(0), G => 
                           first_generate, P => p_vett_0_0_port);
   G_first : GENERAL_G_20 port map( G_in => first_generate, P_in => 
                           p_vett_0_0_port, G_in_prev => Cin, G_out => 
                           g_vett_0_0_port);
   PG_0_1 : PG_block_63 port map( A => A(1), B => B(1), G => g_vett_0_1_port, P
                           => p_vett_0_1_port);
   PG_0_2 : PG_block_62 port map( A => A(2), B => B(2), G => g_vett_0_2_port, P
                           => p_vett_0_2_port);
   PG_0_3 : PG_block_61 port map( A => A(3), B => B(3), G => g_vett_0_3_port, P
                           => p_vett_0_3_port);
   PG_0_4 : PG_block_60 port map( A => A(4), B => B(4), G => g_vett_0_4_port, P
                           => p_vett_0_4_port);
   PG_0_5 : PG_block_59 port map( A => A(5), B => B(5), G => g_vett_0_5_port, P
                           => p_vett_0_5_port);
   PG_0_6 : PG_block_58 port map( A => A(6), B => B(6), G => g_vett_0_6_port, P
                           => p_vett_0_6_port);
   PG_0_7 : PG_block_57 port map( A => A(7), B => B(7), G => g_vett_0_7_port, P
                           => p_vett_0_7_port);
   PG_0_8 : PG_block_56 port map( A => A(8), B => B(8), G => g_vett_0_8_port, P
                           => p_vett_0_8_port);
   PG_0_9 : PG_block_55 port map( A => A(9), B => B(9), G => g_vett_0_9_port, P
                           => p_vett_0_9_port);
   PG_0_10 : PG_block_54 port map( A => A(10), B => B(10), G => 
                           g_vett_0_10_port, P => p_vett_0_10_port);
   PG_0_11 : PG_block_53 port map( A => A(11), B => B(11), G => 
                           g_vett_0_11_port, P => p_vett_0_11_port);
   PG_0_12 : PG_block_52 port map( A => A(12), B => B(12), G => 
                           g_vett_0_12_port, P => p_vett_0_12_port);
   PG_0_13 : PG_block_51 port map( A => A(13), B => B(13), G => 
                           g_vett_0_13_port, P => p_vett_0_13_port);
   PG_0_14 : PG_block_50 port map( A => A(14), B => B(14), G => 
                           g_vett_0_14_port, P => p_vett_0_14_port);
   PG_0_15 : PG_block_49 port map( A => A(15), B => B(15), G => 
                           g_vett_0_15_port, P => p_vett_0_15_port);
   PG_0_16 : PG_block_48 port map( A => A(16), B => B(16), G => 
                           g_vett_0_16_port, P => p_vett_0_16_port);
   PG_0_17 : PG_block_47 port map( A => A(17), B => B(17), G => 
                           g_vett_0_17_port, P => p_vett_0_17_port);
   PG_0_18 : PG_block_46 port map( A => A(18), B => B(18), G => 
                           g_vett_0_18_port, P => p_vett_0_18_port);
   PG_0_19 : PG_block_45 port map( A => A(19), B => B(19), G => 
                           g_vett_0_19_port, P => p_vett_0_19_port);
   PG_0_20 : PG_block_44 port map( A => A(20), B => B(20), G => 
                           g_vett_0_20_port, P => p_vett_0_20_port);
   PG_0_21 : PG_block_43 port map( A => A(21), B => B(21), G => 
                           g_vett_0_21_port, P => p_vett_0_21_port);
   PG_0_22 : PG_block_42 port map( A => A(22), B => B(22), G => 
                           g_vett_0_22_port, P => p_vett_0_22_port);
   PG_0_23 : PG_block_41 port map( A => A(23), B => B(23), G => 
                           g_vett_0_23_port, P => p_vett_0_23_port);
   PG_0_24 : PG_block_40 port map( A => A(24), B => B(24), G => 
                           g_vett_0_24_port, P => p_vett_0_24_port);
   PG_0_25 : PG_block_39 port map( A => A(25), B => B(25), G => 
                           g_vett_0_25_port, P => p_vett_0_25_port);
   PG_0_26 : PG_block_38 port map( A => A(26), B => B(26), G => 
                           g_vett_0_26_port, P => p_vett_0_26_port);
   PG_0_27 : PG_block_37 port map( A => A(27), B => B(27), G => 
                           g_vett_0_27_port, P => p_vett_0_27_port);
   PG_0_28 : PG_block_36 port map( A => A(28), B => B(28), G => 
                           g_vett_0_28_port, P => p_vett_0_28_port);
   PG_0_29 : PG_block_35 port map( A => A(29), B => B(29), G => 
                           g_vett_0_29_port, P => p_vett_0_29_port);
   PG_0_30 : PG_block_34 port map( A => A(30), B => B(30), G => 
                           g_vett_0_30_port, P => p_vett_0_30_port);
   PG_0_31 : PG_block_33 port map( A => A(31), B => B(31), G => 
                           g_vett_0_31_port, P => p_vett_0_31_port);
   G_0_0_0 : GENERAL_G_19 port map( G_in => g_vett_0_1_port, P_in => 
                           p_vett_0_1_port, G_in_prev => g_vett_0_0_port, G_out
                           => g_vett_1_0_port);
   PG_1_0_0 : GENERAL_PG_54 port map( G_in => g_vett_0_3_port, P_in => 
                           p_vett_0_3_port, G_in_prev => g_vett_0_2_port, 
                           P_in_prev => p_vett_0_2_port, G_out => 
                           g_vett_1_1_port, P_out => p_vett_1_1_port);
   G_1_0_0 : GENERAL_G_18 port map( G_in => g_vett_1_1_port, P_in => 
                           p_vett_1_1_port, G_in_prev => g_vett_1_0_port, G_out
                           => Co_1_port);
   PG_2_0_1 : GENERAL_PG_53 port map( G_in => g_vett_0_5_port, P_in => 
                           p_vett_0_5_port, G_in_prev => g_vett_0_4_port, 
                           P_in_prev => p_vett_0_4_port, G_out => 
                           g_vett_1_2_port, P_out => p_vett_1_2_port);
   PG_3_0_1 : GENERAL_PG_52 port map( G_in => g_vett_0_7_port, P_in => 
                           p_vett_0_7_port, G_in_prev => g_vett_0_6_port, 
                           P_in_prev => p_vett_0_6_port, G_out => 
                           g_vett_1_3_port, P_out => p_vett_1_3_port);
   PG_4_0_1 : GENERAL_PG_51 port map( G_in => g_vett_1_3_port, P_in => 
                           p_vett_1_3_port, G_in_prev => g_vett_1_2_port, 
                           P_in_prev => p_vett_1_2_port, G_out => 
                           g_vett_2_1_port, P_out => p_vett_2_1_port);
   PG_2_0_2 : GENERAL_PG_50 port map( G_in => g_vett_0_9_port, P_in => 
                           p_vett_0_9_port, G_in_prev => g_vett_0_8_port, 
                           P_in_prev => p_vett_0_8_port, G_out => 
                           g_vett_1_4_port, P_out => p_vett_1_4_port);
   PG_3_0_2 : GENERAL_PG_49 port map( G_in => g_vett_0_11_port, P_in => 
                           p_vett_0_11_port, G_in_prev => g_vett_0_10_port, 
                           P_in_prev => p_vett_0_10_port, G_out => 
                           g_vett_1_5_port, P_out => p_vett_1_5_port);
   PG_4_0_2 : GENERAL_PG_48 port map( G_in => g_vett_1_5_port, P_in => 
                           p_vett_1_5_port, G_in_prev => g_vett_1_4_port, 
                           P_in_prev => p_vett_1_4_port, G_out => 
                           g_vett_2_2_port, P_out => p_vett_2_2_port);
   PG_2_0_3 : GENERAL_PG_47 port map( G_in => g_vett_0_13_port, P_in => 
                           p_vett_0_13_port, G_in_prev => g_vett_0_12_port, 
                           P_in_prev => p_vett_0_12_port, G_out => 
                           g_vett_1_6_port, P_out => p_vett_1_6_port);
   PG_3_0_3 : GENERAL_PG_46 port map( G_in => g_vett_0_15_port, P_in => 
                           p_vett_0_15_port, G_in_prev => g_vett_0_14_port, 
                           P_in_prev => p_vett_0_14_port, G_out => 
                           g_vett_1_7_port, P_out => p_vett_1_7_port);
   PG_4_0_3 : GENERAL_PG_45 port map( G_in => g_vett_1_7_port, P_in => 
                           p_vett_1_7_port, G_in_prev => g_vett_1_6_port, 
                           P_in_prev => p_vett_1_6_port, G_out => 
                           g_vett_2_3_port, P_out => p_vett_2_3_port);
   PG_2_0_4 : GENERAL_PG_44 port map( G_in => g_vett_0_17_port, P_in => 
                           p_vett_0_17_port, G_in_prev => g_vett_0_16_port, 
                           P_in_prev => p_vett_0_16_port, G_out => 
                           g_vett_1_8_port, P_out => p_vett_1_8_port);
   PG_3_0_4 : GENERAL_PG_43 port map( G_in => g_vett_0_19_port, P_in => 
                           p_vett_0_19_port, G_in_prev => g_vett_0_18_port, 
                           P_in_prev => p_vett_0_18_port, G_out => 
                           g_vett_1_9_port, P_out => p_vett_1_9_port);
   PG_4_0_4 : GENERAL_PG_42 port map( G_in => g_vett_1_9_port, P_in => 
                           p_vett_1_9_port, G_in_prev => g_vett_1_8_port, 
                           P_in_prev => p_vett_1_8_port, G_out => 
                           g_vett_2_4_port, P_out => p_vett_2_4_port);
   PG_2_0_5 : GENERAL_PG_41 port map( G_in => g_vett_0_21_port, P_in => 
                           p_vett_0_21_port, G_in_prev => g_vett_0_20_port, 
                           P_in_prev => p_vett_0_20_port, G_out => 
                           g_vett_1_10_port, P_out => p_vett_1_10_port);
   PG_3_0_5 : GENERAL_PG_40 port map( G_in => g_vett_0_23_port, P_in => 
                           p_vett_0_23_port, G_in_prev => g_vett_0_22_port, 
                           P_in_prev => p_vett_0_22_port, G_out => 
                           g_vett_1_11_port, P_out => p_vett_1_11_port);
   PG_4_0_5 : GENERAL_PG_39 port map( G_in => g_vett_1_11_port, P_in => 
                           p_vett_1_11_port, G_in_prev => g_vett_1_10_port, 
                           P_in_prev => p_vett_1_10_port, G_out => 
                           g_vett_2_5_port, P_out => p_vett_2_5_port);
   PG_2_0_6 : GENERAL_PG_38 port map( G_in => g_vett_0_25_port, P_in => 
                           p_vett_0_25_port, G_in_prev => g_vett_0_24_port, 
                           P_in_prev => p_vett_0_24_port, G_out => 
                           g_vett_1_12_port, P_out => p_vett_1_12_port);
   PG_3_0_6 : GENERAL_PG_37 port map( G_in => g_vett_0_27_port, P_in => 
                           p_vett_0_27_port, G_in_prev => g_vett_0_26_port, 
                           P_in_prev => p_vett_0_26_port, G_out => 
                           g_vett_1_13_port, P_out => p_vett_1_13_port);
   PG_4_0_6 : GENERAL_PG_36 port map( G_in => g_vett_1_13_port, P_in => 
                           p_vett_1_13_port, G_in_prev => g_vett_1_12_port, 
                           P_in_prev => p_vett_1_12_port, G_out => 
                           g_vett_2_6_port, P_out => p_vett_2_6_port);
   PG_2_0_7 : GENERAL_PG_35 port map( G_in => g_vett_0_29_port, P_in => 
                           p_vett_0_29_port, G_in_prev => g_vett_0_28_port, 
                           P_in_prev => p_vett_0_28_port, G_out => 
                           g_vett_1_14_port, P_out => p_vett_1_14_port);
   PG_3_0_7 : GENERAL_PG_34 port map( G_in => g_vett_0_31_port, P_in => 
                           p_vett_0_31_port, G_in_prev => g_vett_0_30_port, 
                           P_in_prev => p_vett_0_30_port, G_out => 
                           g_vett_1_15_port, P_out => p_vett_1_15_port);
   PG_4_0_7 : GENERAL_PG_33 port map( G_in => g_vett_1_15_port, P_in => 
                           p_vett_1_15_port, G_in_prev => g_vett_1_14_port, 
                           P_in_prev => p_vett_1_14_port, G_out => 
                           g_vett_2_7_port, P_out => p_vett_2_7_port);
   G_2_1_0 : GENERAL_G_17 port map( G_in => g_vett_2_1_port, P_in => 
                           p_vett_2_1_port, G_in_prev => Co_1_port, G_out => 
                           Co_2_port);
   PG_5_1_0 : GENERAL_PG_32 port map( G_in => g_vett_2_3_port, P_in => 
                           p_vett_2_3_port, G_in_prev => g_vett_2_2_port, 
                           P_in_prev => p_vett_2_2_port, G_out => 
                           g_vett_3_1_port, P_out => p_vett_3_1_port);
   G_3_1_0 : GENERAL_G_16 port map( G_in => g_vett_2_2_port, P_in => 
                           p_vett_2_2_port, G_in_prev => Co_2_port, G_out => 
                           Co_3_port);
   G_4_1_0 : GENERAL_G_15 port map( G_in => g_vett_3_1_port, P_in => 
                           p_vett_3_1_port, G_in_prev => Co_2_port, G_out => 
                           Co_4_port);
   PG_6_1_1 : GENERAL_PG_31 port map( G_in => g_vett_2_5_port, P_in => 
                           p_vett_2_5_port, G_in_prev => g_vett_2_4_port, 
                           P_in_prev => p_vett_2_4_port, G_out => 
                           g_vett_3_2_port, P_out => p_vett_3_2_port);
   PG_7_1_1 : GENERAL_PG_30 port map( G_in => g_vett_2_7_port, P_in => 
                           p_vett_2_7_port, G_in_prev => g_vett_2_6_port, 
                           P_in_prev => p_vett_2_6_port, G_out => 
                           g_vett_3_3_port, P_out => p_vett_3_3_port);
   PG_8_1_1 : GENERAL_PG_29 port map( G_in => g_vett_2_6_port, P_in => 
                           p_vett_2_6_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_2_port, P_out => p_vett_4_2_port);
   PG_9_1_1 : GENERAL_PG_28 port map( G_in => g_vett_3_3_port, P_in => 
                           p_vett_3_3_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_3_port, P_out => p_vett_4_3_port);
   G_5_2_0 : GENERAL_G_14 port map( G_in => g_vett_2_4_port, P_in => 
                           p_vett_2_4_port, G_in_prev => Co_4_port, G_out => 
                           Co_5_port);
   G_6_2_1 : GENERAL_G_13 port map( G_in => g_vett_3_2_port, P_in => 
                           p_vett_3_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_6_port);
   G_7_2_2 : GENERAL_G_12 port map( G_in => g_vett_4_2_port, P_in => 
                           p_vett_4_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_7_port);
   G_8_2_3 : GENERAL_G_11 port map( G_in => g_vett_4_3_port, P_in => 
                           p_vett_4_3_port, G_in_prev => Co_4_port, G_out => 
                           n_1115);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity SUMGEN_NBIT32_NBLOCKS8_3 is

   port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
         std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
         std_logic_vector (31 downto 0));

end SUMGEN_NBIT32_NBLOCKS8_3;

architecture SYN_STRUCTURAL of SUMGEN_NBIT32_NBLOCKS8_3 is

   component CSblock_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122 : std_logic;

begin
   
   block_i_0 : CSblock_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), cin => cin_vect(0), Y(3) => 
                           SUM(3), Y(2) => SUM(2), Y(1) => SUM(1), Y(0) => 
                           SUM(0), Co => n_1116);
   block_i_1 : CSblock_NBIT4_23 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), cin => cin_vect(1), Y(3) => 
                           SUM(7), Y(2) => SUM(6), Y(1) => SUM(5), Y(0) => 
                           SUM(4), Co => n_1117);
   block_i_2 : CSblock_NBIT4_22 port map( A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), cin => cin_vect(2), Y(3)
                           => SUM(11), Y(2) => SUM(10), Y(1) => SUM(9), Y(0) =>
                           SUM(8), Co => n_1118);
   block_i_3 : CSblock_NBIT4_21 port map( A(3) => A(15), A(2) => A(14), A(1) =>
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), cin => cin_vect(3), 
                           Y(3) => SUM(15), Y(2) => SUM(14), Y(1) => SUM(13), 
                           Y(0) => SUM(12), Co => n_1119);
   block_i_4 : CSblock_NBIT4_20 port map( A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), cin => cin_vect(4), 
                           Y(3) => SUM(19), Y(2) => SUM(18), Y(1) => SUM(17), 
                           Y(0) => SUM(16), Co => n_1120);
   block_i_5 : CSblock_NBIT4_19 port map( A(3) => A(23), A(2) => A(22), A(1) =>
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), cin => cin_vect(5), 
                           Y(3) => SUM(23), Y(2) => SUM(22), Y(1) => SUM(21), 
                           Y(0) => SUM(20), Co => n_1121);
   block_i_6 : CSblock_NBIT4_18 port map( A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), cin => cin_vect(6), 
                           Y(3) => SUM(27), Y(2) => SUM(26), Y(1) => SUM(25), 
                           Y(0) => SUM(24), Co => n_1122);
   block_i_7 : CSblock_NBIT4_17 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), cin => cin_vect(7), 
                           Y(3) => SUM(31), Y(2) => SUM(30), Y(1) => SUM(29), 
                           Y(0) => SUM(28), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 is

   component GENERAL_G_21
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_22
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_23
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_24
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_55
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_56
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_57
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_58
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_25
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_26
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_59
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_27
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_60
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_61
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_62
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_63
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_64
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_65
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_66
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_67
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_68
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_69
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_70
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_71
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_72
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_73
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_74
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_75
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_76
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_77
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_78
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_79
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_80
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_28
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_81
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_29
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_65
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_66
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_67
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_68
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_69
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_70
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_71
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_72
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_73
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_74
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_75
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_76
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_77
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_78
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_79
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_80
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_81
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_82
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_83
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_84
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_85
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_86
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_87
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_88
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_89
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_90
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_91
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_92
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_93
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_94
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_95
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component GENERAL_G_30
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_96
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, first_generate, p_vett_4_3_port, p_vett_4_2_port, 
      p_vett_3_3_port, p_vett_3_2_port, p_vett_3_1_port, p_vett_2_7_port, 
      p_vett_2_6_port, p_vett_2_5_port, p_vett_2_4_port, p_vett_2_3_port, 
      p_vett_2_2_port, p_vett_2_1_port, p_vett_1_15_port, p_vett_1_14_port, 
      p_vett_1_13_port, p_vett_1_12_port, p_vett_1_11_port, p_vett_1_10_port, 
      p_vett_1_9_port, p_vett_1_8_port, p_vett_1_7_port, p_vett_1_6_port, 
      p_vett_1_5_port, p_vett_1_4_port, p_vett_1_3_port, p_vett_1_2_port, 
      p_vett_1_1_port, p_vett_0_31_port, p_vett_0_30_port, p_vett_0_29_port, 
      p_vett_0_28_port, p_vett_0_27_port, p_vett_0_26_port, p_vett_0_25_port, 
      p_vett_0_24_port, p_vett_0_23_port, p_vett_0_22_port, p_vett_0_21_port, 
      p_vett_0_20_port, p_vett_0_19_port, p_vett_0_18_port, p_vett_0_17_port, 
      p_vett_0_16_port, p_vett_0_15_port, p_vett_0_14_port, p_vett_0_13_port, 
      p_vett_0_12_port, p_vett_0_11_port, p_vett_0_10_port, p_vett_0_9_port, 
      p_vett_0_8_port, p_vett_0_7_port, p_vett_0_6_port, p_vett_0_5_port, 
      p_vett_0_4_port, p_vett_0_3_port, p_vett_0_2_port, p_vett_0_1_port, 
      p_vett_0_0_port, g_vett_4_3_port, g_vett_4_2_port, g_vett_3_3_port, 
      g_vett_3_2_port, g_vett_3_1_port, g_vett_2_7_port, g_vett_2_6_port, 
      g_vett_2_5_port, g_vett_2_4_port, g_vett_2_3_port, g_vett_2_2_port, 
      g_vett_2_1_port, g_vett_1_15_port, g_vett_1_14_port, g_vett_1_13_port, 
      g_vett_1_12_port, g_vett_1_11_port, g_vett_1_10_port, g_vett_1_9_port, 
      g_vett_1_8_port, g_vett_1_7_port, g_vett_1_6_port, g_vett_1_5_port, 
      g_vett_1_4_port, g_vett_1_3_port, g_vett_1_2_port, g_vett_1_1_port, 
      g_vett_1_0_port, g_vett_0_31_port, g_vett_0_30_port, g_vett_0_29_port, 
      g_vett_0_28_port, g_vett_0_27_port, g_vett_0_26_port, g_vett_0_25_port, 
      g_vett_0_24_port, g_vett_0_23_port, g_vett_0_22_port, g_vett_0_21_port, 
      g_vett_0_20_port, g_vett_0_19_port, g_vett_0_18_port, g_vett_0_17_port, 
      g_vett_0_16_port, g_vett_0_15_port, g_vett_0_14_port, g_vett_0_13_port, 
      g_vett_0_12_port, g_vett_0_11_port, g_vett_0_10_port, g_vett_0_9_port, 
      g_vett_0_8_port, g_vett_0_7_port, g_vett_0_6_port, g_vett_0_5_port, 
      g_vett_0_4_port, g_vett_0_3_port, g_vett_0_2_port, g_vett_0_1_port, 
      g_vett_0_0_port, n_1123 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Cin );
   
   PGblock_first : PG_block_96 port map( A => A(0), B => B(0), G => 
                           first_generate, P => p_vett_0_0_port);
   G_first : GENERAL_G_30 port map( G_in => first_generate, P_in => 
                           p_vett_0_0_port, G_in_prev => Cin, G_out => 
                           g_vett_0_0_port);
   PG_0_1 : PG_block_95 port map( A => A(1), B => B(1), G => g_vett_0_1_port, P
                           => p_vett_0_1_port);
   PG_0_2 : PG_block_94 port map( A => A(2), B => B(2), G => g_vett_0_2_port, P
                           => p_vett_0_2_port);
   PG_0_3 : PG_block_93 port map( A => A(3), B => B(3), G => g_vett_0_3_port, P
                           => p_vett_0_3_port);
   PG_0_4 : PG_block_92 port map( A => A(4), B => B(4), G => g_vett_0_4_port, P
                           => p_vett_0_4_port);
   PG_0_5 : PG_block_91 port map( A => A(5), B => B(5), G => g_vett_0_5_port, P
                           => p_vett_0_5_port);
   PG_0_6 : PG_block_90 port map( A => A(6), B => B(6), G => g_vett_0_6_port, P
                           => p_vett_0_6_port);
   PG_0_7 : PG_block_89 port map( A => A(7), B => B(7), G => g_vett_0_7_port, P
                           => p_vett_0_7_port);
   PG_0_8 : PG_block_88 port map( A => A(8), B => B(8), G => g_vett_0_8_port, P
                           => p_vett_0_8_port);
   PG_0_9 : PG_block_87 port map( A => A(9), B => B(9), G => g_vett_0_9_port, P
                           => p_vett_0_9_port);
   PG_0_10 : PG_block_86 port map( A => A(10), B => B(10), G => 
                           g_vett_0_10_port, P => p_vett_0_10_port);
   PG_0_11 : PG_block_85 port map( A => A(11), B => B(11), G => 
                           g_vett_0_11_port, P => p_vett_0_11_port);
   PG_0_12 : PG_block_84 port map( A => A(12), B => B(12), G => 
                           g_vett_0_12_port, P => p_vett_0_12_port);
   PG_0_13 : PG_block_83 port map( A => A(13), B => B(13), G => 
                           g_vett_0_13_port, P => p_vett_0_13_port);
   PG_0_14 : PG_block_82 port map( A => A(14), B => B(14), G => 
                           g_vett_0_14_port, P => p_vett_0_14_port);
   PG_0_15 : PG_block_81 port map( A => A(15), B => B(15), G => 
                           g_vett_0_15_port, P => p_vett_0_15_port);
   PG_0_16 : PG_block_80 port map( A => A(16), B => B(16), G => 
                           g_vett_0_16_port, P => p_vett_0_16_port);
   PG_0_17 : PG_block_79 port map( A => A(17), B => B(17), G => 
                           g_vett_0_17_port, P => p_vett_0_17_port);
   PG_0_18 : PG_block_78 port map( A => A(18), B => B(18), G => 
                           g_vett_0_18_port, P => p_vett_0_18_port);
   PG_0_19 : PG_block_77 port map( A => A(19), B => B(19), G => 
                           g_vett_0_19_port, P => p_vett_0_19_port);
   PG_0_20 : PG_block_76 port map( A => A(20), B => B(20), G => 
                           g_vett_0_20_port, P => p_vett_0_20_port);
   PG_0_21 : PG_block_75 port map( A => A(21), B => B(21), G => 
                           g_vett_0_21_port, P => p_vett_0_21_port);
   PG_0_22 : PG_block_74 port map( A => A(22), B => B(22), G => 
                           g_vett_0_22_port, P => p_vett_0_22_port);
   PG_0_23 : PG_block_73 port map( A => A(23), B => B(23), G => 
                           g_vett_0_23_port, P => p_vett_0_23_port);
   PG_0_24 : PG_block_72 port map( A => A(24), B => B(24), G => 
                           g_vett_0_24_port, P => p_vett_0_24_port);
   PG_0_25 : PG_block_71 port map( A => A(25), B => B(25), G => 
                           g_vett_0_25_port, P => p_vett_0_25_port);
   PG_0_26 : PG_block_70 port map( A => A(26), B => B(26), G => 
                           g_vett_0_26_port, P => p_vett_0_26_port);
   PG_0_27 : PG_block_69 port map( A => A(27), B => B(27), G => 
                           g_vett_0_27_port, P => p_vett_0_27_port);
   PG_0_28 : PG_block_68 port map( A => A(28), B => B(28), G => 
                           g_vett_0_28_port, P => p_vett_0_28_port);
   PG_0_29 : PG_block_67 port map( A => A(29), B => B(29), G => 
                           g_vett_0_29_port, P => p_vett_0_29_port);
   PG_0_30 : PG_block_66 port map( A => A(30), B => B(30), G => 
                           g_vett_0_30_port, P => p_vett_0_30_port);
   PG_0_31 : PG_block_65 port map( A => A(31), B => B(31), G => 
                           g_vett_0_31_port, P => p_vett_0_31_port);
   G_0_0_0 : GENERAL_G_29 port map( G_in => g_vett_0_1_port, P_in => 
                           p_vett_0_1_port, G_in_prev => g_vett_0_0_port, G_out
                           => g_vett_1_0_port);
   PG_1_0_0 : GENERAL_PG_81 port map( G_in => g_vett_0_3_port, P_in => 
                           p_vett_0_3_port, G_in_prev => g_vett_0_2_port, 
                           P_in_prev => p_vett_0_2_port, G_out => 
                           g_vett_1_1_port, P_out => p_vett_1_1_port);
   G_1_0_0 : GENERAL_G_28 port map( G_in => g_vett_1_1_port, P_in => 
                           p_vett_1_1_port, G_in_prev => g_vett_1_0_port, G_out
                           => Co_1_port);
   PG_2_0_1 : GENERAL_PG_80 port map( G_in => g_vett_0_5_port, P_in => 
                           p_vett_0_5_port, G_in_prev => g_vett_0_4_port, 
                           P_in_prev => p_vett_0_4_port, G_out => 
                           g_vett_1_2_port, P_out => p_vett_1_2_port);
   PG_3_0_1 : GENERAL_PG_79 port map( G_in => g_vett_0_7_port, P_in => 
                           p_vett_0_7_port, G_in_prev => g_vett_0_6_port, 
                           P_in_prev => p_vett_0_6_port, G_out => 
                           g_vett_1_3_port, P_out => p_vett_1_3_port);
   PG_4_0_1 : GENERAL_PG_78 port map( G_in => g_vett_1_3_port, P_in => 
                           p_vett_1_3_port, G_in_prev => g_vett_1_2_port, 
                           P_in_prev => p_vett_1_2_port, G_out => 
                           g_vett_2_1_port, P_out => p_vett_2_1_port);
   PG_2_0_2 : GENERAL_PG_77 port map( G_in => g_vett_0_9_port, P_in => 
                           p_vett_0_9_port, G_in_prev => g_vett_0_8_port, 
                           P_in_prev => p_vett_0_8_port, G_out => 
                           g_vett_1_4_port, P_out => p_vett_1_4_port);
   PG_3_0_2 : GENERAL_PG_76 port map( G_in => g_vett_0_11_port, P_in => 
                           p_vett_0_11_port, G_in_prev => g_vett_0_10_port, 
                           P_in_prev => p_vett_0_10_port, G_out => 
                           g_vett_1_5_port, P_out => p_vett_1_5_port);
   PG_4_0_2 : GENERAL_PG_75 port map( G_in => g_vett_1_5_port, P_in => 
                           p_vett_1_5_port, G_in_prev => g_vett_1_4_port, 
                           P_in_prev => p_vett_1_4_port, G_out => 
                           g_vett_2_2_port, P_out => p_vett_2_2_port);
   PG_2_0_3 : GENERAL_PG_74 port map( G_in => g_vett_0_13_port, P_in => 
                           p_vett_0_13_port, G_in_prev => g_vett_0_12_port, 
                           P_in_prev => p_vett_0_12_port, G_out => 
                           g_vett_1_6_port, P_out => p_vett_1_6_port);
   PG_3_0_3 : GENERAL_PG_73 port map( G_in => g_vett_0_15_port, P_in => 
                           p_vett_0_15_port, G_in_prev => g_vett_0_14_port, 
                           P_in_prev => p_vett_0_14_port, G_out => 
                           g_vett_1_7_port, P_out => p_vett_1_7_port);
   PG_4_0_3 : GENERAL_PG_72 port map( G_in => g_vett_1_7_port, P_in => 
                           p_vett_1_7_port, G_in_prev => g_vett_1_6_port, 
                           P_in_prev => p_vett_1_6_port, G_out => 
                           g_vett_2_3_port, P_out => p_vett_2_3_port);
   PG_2_0_4 : GENERAL_PG_71 port map( G_in => g_vett_0_17_port, P_in => 
                           p_vett_0_17_port, G_in_prev => g_vett_0_16_port, 
                           P_in_prev => p_vett_0_16_port, G_out => 
                           g_vett_1_8_port, P_out => p_vett_1_8_port);
   PG_3_0_4 : GENERAL_PG_70 port map( G_in => g_vett_0_19_port, P_in => 
                           p_vett_0_19_port, G_in_prev => g_vett_0_18_port, 
                           P_in_prev => p_vett_0_18_port, G_out => 
                           g_vett_1_9_port, P_out => p_vett_1_9_port);
   PG_4_0_4 : GENERAL_PG_69 port map( G_in => g_vett_1_9_port, P_in => 
                           p_vett_1_9_port, G_in_prev => g_vett_1_8_port, 
                           P_in_prev => p_vett_1_8_port, G_out => 
                           g_vett_2_4_port, P_out => p_vett_2_4_port);
   PG_2_0_5 : GENERAL_PG_68 port map( G_in => g_vett_0_21_port, P_in => 
                           p_vett_0_21_port, G_in_prev => g_vett_0_20_port, 
                           P_in_prev => p_vett_0_20_port, G_out => 
                           g_vett_1_10_port, P_out => p_vett_1_10_port);
   PG_3_0_5 : GENERAL_PG_67 port map( G_in => g_vett_0_23_port, P_in => 
                           p_vett_0_23_port, G_in_prev => g_vett_0_22_port, 
                           P_in_prev => p_vett_0_22_port, G_out => 
                           g_vett_1_11_port, P_out => p_vett_1_11_port);
   PG_4_0_5 : GENERAL_PG_66 port map( G_in => g_vett_1_11_port, P_in => 
                           p_vett_1_11_port, G_in_prev => g_vett_1_10_port, 
                           P_in_prev => p_vett_1_10_port, G_out => 
                           g_vett_2_5_port, P_out => p_vett_2_5_port);
   PG_2_0_6 : GENERAL_PG_65 port map( G_in => g_vett_0_25_port, P_in => 
                           p_vett_0_25_port, G_in_prev => g_vett_0_24_port, 
                           P_in_prev => p_vett_0_24_port, G_out => 
                           g_vett_1_12_port, P_out => p_vett_1_12_port);
   PG_3_0_6 : GENERAL_PG_64 port map( G_in => g_vett_0_27_port, P_in => 
                           p_vett_0_27_port, G_in_prev => g_vett_0_26_port, 
                           P_in_prev => p_vett_0_26_port, G_out => 
                           g_vett_1_13_port, P_out => p_vett_1_13_port);
   PG_4_0_6 : GENERAL_PG_63 port map( G_in => g_vett_1_13_port, P_in => 
                           p_vett_1_13_port, G_in_prev => g_vett_1_12_port, 
                           P_in_prev => p_vett_1_12_port, G_out => 
                           g_vett_2_6_port, P_out => p_vett_2_6_port);
   PG_2_0_7 : GENERAL_PG_62 port map( G_in => g_vett_0_29_port, P_in => 
                           p_vett_0_29_port, G_in_prev => g_vett_0_28_port, 
                           P_in_prev => p_vett_0_28_port, G_out => 
                           g_vett_1_14_port, P_out => p_vett_1_14_port);
   PG_3_0_7 : GENERAL_PG_61 port map( G_in => g_vett_0_31_port, P_in => 
                           p_vett_0_31_port, G_in_prev => g_vett_0_30_port, 
                           P_in_prev => p_vett_0_30_port, G_out => 
                           g_vett_1_15_port, P_out => p_vett_1_15_port);
   PG_4_0_7 : GENERAL_PG_60 port map( G_in => g_vett_1_15_port, P_in => 
                           p_vett_1_15_port, G_in_prev => g_vett_1_14_port, 
                           P_in_prev => p_vett_1_14_port, G_out => 
                           g_vett_2_7_port, P_out => p_vett_2_7_port);
   G_2_1_0 : GENERAL_G_27 port map( G_in => g_vett_2_1_port, P_in => 
                           p_vett_2_1_port, G_in_prev => Co_1_port, G_out => 
                           Co_2_port);
   PG_5_1_0 : GENERAL_PG_59 port map( G_in => g_vett_2_3_port, P_in => 
                           p_vett_2_3_port, G_in_prev => g_vett_2_2_port, 
                           P_in_prev => p_vett_2_2_port, G_out => 
                           g_vett_3_1_port, P_out => p_vett_3_1_port);
   G_3_1_0 : GENERAL_G_26 port map( G_in => g_vett_2_2_port, P_in => 
                           p_vett_2_2_port, G_in_prev => Co_2_port, G_out => 
                           Co_3_port);
   G_4_1_0 : GENERAL_G_25 port map( G_in => g_vett_3_1_port, P_in => 
                           p_vett_3_1_port, G_in_prev => Co_2_port, G_out => 
                           Co_4_port);
   PG_6_1_1 : GENERAL_PG_58 port map( G_in => g_vett_2_5_port, P_in => 
                           p_vett_2_5_port, G_in_prev => g_vett_2_4_port, 
                           P_in_prev => p_vett_2_4_port, G_out => 
                           g_vett_3_2_port, P_out => p_vett_3_2_port);
   PG_7_1_1 : GENERAL_PG_57 port map( G_in => g_vett_2_7_port, P_in => 
                           p_vett_2_7_port, G_in_prev => g_vett_2_6_port, 
                           P_in_prev => p_vett_2_6_port, G_out => 
                           g_vett_3_3_port, P_out => p_vett_3_3_port);
   PG_8_1_1 : GENERAL_PG_56 port map( G_in => g_vett_2_6_port, P_in => 
                           p_vett_2_6_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_2_port, P_out => p_vett_4_2_port);
   PG_9_1_1 : GENERAL_PG_55 port map( G_in => g_vett_3_3_port, P_in => 
                           p_vett_3_3_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_3_port, P_out => p_vett_4_3_port);
   G_5_2_0 : GENERAL_G_24 port map( G_in => g_vett_2_4_port, P_in => 
                           p_vett_2_4_port, G_in_prev => Co_4_port, G_out => 
                           Co_5_port);
   G_6_2_1 : GENERAL_G_23 port map( G_in => g_vett_3_2_port, P_in => 
                           p_vett_3_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_6_port);
   G_7_2_2 : GENERAL_G_22 port map( G_in => g_vett_4_2_port, P_in => 
                           p_vett_4_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_7_port);
   G_8_2_3 : GENERAL_G_21 port map( G_in => g_vett_4_3_port, P_in => 
                           p_vett_4_3_port, G_in_prev => Co_4_port, G_out => 
                           n_1123);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity mux11to1_nbit32 is

   port( A, B, C, D, E, F, H : in std_logic_vector (31 downto 0);  sel : in 
         std_logic_vector (3 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux11to1_nbit32;

architecture SYN_beh of mux11to1_nbit32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n107, n108,
      net52587, net56040, net56038, net56036, net56046, net56044, net56042, 
      net56052, net56050, net56048, net56058, net56056, net56054, net56064, 
      net56062, net56060, net56070, net56068, net56066, net56076, net56074, 
      net56072, n11, n105, n10, n109, n110, n111, n112, n113, n114, n115, n116,
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153 : std_logic;

begin
   
   U110 : NAND3_X1 port map( A1 => n4, A2 => n5, A3 => n6, ZN => Y(9));
   U111 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => Y(8));
   U113 : NAND3_X1 port map( A1 => n20, A2 => n21, A3 => n22, ZN => Y(6));
   U115 : NAND3_X1 port map( A1 => n26, A2 => n27, A3 => n28, ZN => Y(4));
   U116 : NAND3_X1 port map( A1 => n29, A2 => n30, A3 => n31, ZN => Y(3));
   U118 : NAND3_X1 port map( A1 => n35, A2 => n36, A3 => n37, ZN => Y(30));
   U119 : NAND3_X1 port map( A1 => n40, A2 => n39, A3 => n38, ZN => Y(2));
   U120 : NAND3_X1 port map( A1 => n41, A2 => n42, A3 => n43, ZN => Y(29));
   U121 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => n46, ZN => Y(28));
   U122 : NAND3_X1 port map( A1 => n47, A2 => n48, A3 => n49, ZN => Y(27));
   U123 : NAND3_X1 port map( A1 => n50, A2 => n51, A3 => n52, ZN => Y(26));
   U124 : NAND3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => Y(25));
   U125 : NAND3_X1 port map( A1 => n56, A2 => n57, A3 => n58, ZN => Y(24));
   U126 : NAND3_X1 port map( A1 => n59, A2 => n60, A3 => n61, ZN => Y(23));
   U127 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => Y(22));
   U128 : NAND3_X1 port map( A1 => n65, A2 => n66, A3 => n67, ZN => Y(21));
   U129 : NAND3_X1 port map( A1 => n68, A2 => n69, A3 => n70, ZN => Y(20));
   U130 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => Y(1));
   U131 : NAND3_X1 port map( A1 => n74, A2 => n75, A3 => n76, ZN => Y(19));
   U132 : NAND3_X1 port map( A1 => n77, A2 => n78, A3 => n79, ZN => Y(18));
   U133 : NAND3_X1 port map( A1 => n82, A2 => n81, A3 => n80, ZN => Y(17));
   U134 : NAND3_X1 port map( A1 => n83, A2 => n84, A3 => n85, ZN => Y(16));
   U135 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n88, ZN => Y(15));
   U136 : NAND3_X1 port map( A1 => n89, A2 => n90, A3 => n91, ZN => Y(14));
   U137 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n94, ZN => Y(13));
   U140 : NAND3_X1 port map( A1 => n101, A2 => n102, A3 => n103, ZN => Y(10));
   U2 : BUF_X1 port map( A => n9, Z => net56048);
   U3 : BUF_X1 port map( A => n9, Z => net56050);
   U4 : AND2_X1 port map( A1 => n131, A2 => n132, ZN => n126);
   U5 : AND2_X1 port map( A1 => n34, A2 => n33, ZN => n109);
   U6 : AND2_X1 port map( A1 => n95, A2 => n96, ZN => n110);
   U7 : AND2_X1 port map( A1 => n98, A2 => n99, ZN => n111);
   U8 : AND2_X1 port map( A1 => n17, A2 => n18, ZN => n112);
   U9 : INV_X1 port map( A => n104, ZN => n115);
   U10 : AND2_X1 port map( A1 => n23, A2 => n24, ZN => n113);
   U11 : NOR2_X1 port map( A1 => n116, A2 => n115, ZN => n114);
   U12 : NAND3_X1 port map( A1 => n140, A2 => n141, A3 => n142, ZN => n116);
   U13 : AOI22_X1 port map( A1 => E(4), A2 => net56070, B1 => C(4), B2 => 
                           net56076, ZN => n26);
   U14 : NAND2_X1 port map( A1 => A(18), A2 => net56036, ZN => n117);
   U15 : NAND2_X1 port map( A1 => B(18), A2 => net56042, ZN => n118);
   U16 : NAND2_X1 port map( A1 => F(18), A2 => net56048, ZN => n119);
   U17 : AND3_X1 port map( A1 => n117, A2 => n118, A3 => n119, ZN => n79);
   U18 : NAND2_X1 port map( A1 => A(6), A2 => net56040, ZN => n120);
   U19 : NAND2_X1 port map( A1 => B(6), A2 => net56046, ZN => n121);
   U20 : NAND2_X1 port map( A1 => F(6), A2 => net56052, ZN => n122);
   U21 : AND3_X1 port map( A1 => n120, A2 => n121, A3 => n122, ZN => n22);
   U22 : NAND2_X1 port map( A1 => A(1), A2 => net56036, ZN => n123);
   U23 : NAND2_X1 port map( A1 => B(1), A2 => net56042, ZN => n124);
   U24 : NAND2_X1 port map( A1 => F(1), A2 => net56048, ZN => n125);
   U25 : AND3_X1 port map( A1 => n123, A2 => n124, A3 => n125, ZN => n73);
   U26 : AND2_X1 port map( A1 => n133, A2 => n126, ZN => n97);
   U27 : NAND2_X1 port map( A1 => n19, A2 => n112, ZN => Y(7));
   U28 : NAND2_X1 port map( A1 => n97, A2 => n110, ZN => Y(12));
   U29 : NAND2_X1 port map( A1 => A(4), A2 => net56040, ZN => n127);
   U30 : NAND2_X1 port map( A1 => B(4), A2 => net56046, ZN => n128);
   U31 : NAND2_X1 port map( A1 => F(4), A2 => net56052, ZN => n129);
   U32 : AND3_X1 port map( A1 => n127, A2 => n128, A3 => n129, ZN => n28);
   U33 : BUF_X1 port map( A => n9, Z => net56052);
   U34 : AND2_X1 port map( A1 => n134, A2 => n135, ZN => n130);
   U35 : AND2_X1 port map( A1 => n136, A2 => n130, ZN => n100);
   U36 : NAND2_X1 port map( A1 => n100, A2 => n111, ZN => Y(11));
   U37 : NAND2_X1 port map( A1 => A(12), A2 => net56036, ZN => n131);
   U38 : NAND2_X1 port map( A1 => B(12), A2 => net56042, ZN => n132);
   U39 : NAND2_X1 port map( A1 => F(12), A2 => net56048, ZN => n133);
   U40 : NAND2_X1 port map( A1 => A(11), A2 => net56036, ZN => n134);
   U41 : NAND2_X1 port map( A1 => B(11), A2 => net56042, ZN => n135);
   U42 : NAND2_X1 port map( A1 => F(11), A2 => net56048, ZN => n136);
   U43 : NAND2_X1 port map( A1 => A(7), A2 => net56040, ZN => n137);
   U44 : NAND2_X1 port map( A1 => B(7), A2 => net56046, ZN => n138);
   U45 : NAND2_X1 port map( A1 => F(7), A2 => net56052, ZN => n139);
   U46 : AND3_X1 port map( A1 => n137, A2 => n138, A3 => n139, ZN => n19);
   U47 : NAND2_X1 port map( A1 => A(0), A2 => net56036, ZN => n140);
   U48 : NAND2_X1 port map( A1 => B(0), A2 => net56042, ZN => n141);
   U49 : NAND2_X1 port map( A1 => F(0), A2 => net56048, ZN => n142);
   U50 : NAND2_X1 port map( A1 => n25, A2 => n113, ZN => Y(5));
   U51 : NAND2_X1 port map( A1 => A(9), A2 => net56040, ZN => n143);
   U52 : NAND2_X1 port map( A1 => B(9), A2 => net56046, ZN => n144);
   U53 : NAND2_X1 port map( A1 => F(9), A2 => net56052, ZN => n145);
   U54 : AND3_X1 port map( A1 => n143, A2 => n144, A3 => n145, ZN => n6);
   U55 : NAND2_X1 port map( A1 => A(2), A2 => net56038, ZN => n146);
   U56 : NAND2_X1 port map( A1 => B(2), A2 => net56044, ZN => n147);
   U57 : NAND2_X1 port map( A1 => F(2), A2 => net56050, ZN => n148);
   U58 : AND3_X1 port map( A1 => n148, A2 => n147, A3 => n146, ZN => n40);
   U59 : AOI22_X1 port map( A1 => D(0), A2 => net56054, B1 => H(0), B2 => 
                           net56060, ZN => n105);
   U60 : NAND2_X1 port map( A1 => n105, A2 => n114, ZN => Y(0));
   U61 : BUF_X1 port map( A => n11, Z => net56060);
   U62 : BUF_X1 port map( A => n10, Z => net56054);
   U63 : AND3_X1 port map( A1 => sel(1), A2 => sel(0), A3 => n107, ZN => n11);
   U64 : BUF_X1 port map( A => n11, Z => net56062);
   U65 : BUF_X1 port map( A => n11, Z => net56064);
   U66 : AND3_X1 port map( A1 => sel(0), A2 => n108, A3 => sel(1), ZN => n10);
   U67 : BUF_X1 port map( A => n10, Z => net56056);
   U68 : BUF_X1 port map( A => n10, Z => net56058);
   U69 : AND3_X1 port map( A1 => n108, A2 => net52587, A3 => sel(1), ZN => n13)
                           ;
   U70 : INV_X1 port map( A => sel(1), ZN => n149);
   U71 : AND3_X1 port map( A1 => net52587, A2 => n149, A3 => n107, ZN => n12);
   U72 : AND3_X1 port map( A1 => sel(0), A2 => n149, A3 => n107, ZN => n9);
   U73 : AND3_X1 port map( A1 => net52587, A2 => n149, A3 => n108, ZN => n7);
   U74 : AND3_X1 port map( A1 => n108, A2 => n149, A3 => sel(0), ZN => n8);
   U75 : NAND2_X1 port map( A1 => n32, A2 => n109, ZN => Y(31));
   U76 : NAND2_X1 port map( A1 => A(5), A2 => net56040, ZN => n150);
   U77 : NAND2_X1 port map( A1 => B(5), A2 => net56046, ZN => n151);
   U78 : NAND2_X1 port map( A1 => F(5), A2 => net56052, ZN => n152);
   U79 : AND3_X1 port map( A1 => n150, A2 => n151, A3 => n152, ZN => n25);
   U80 : BUF_X1 port map( A => n12, Z => net56066);
   U81 : BUF_X1 port map( A => n12, Z => net56068);
   U82 : BUF_X1 port map( A => n7, Z => net56038);
   U83 : BUF_X1 port map( A => n7, Z => net56036);
   U84 : BUF_X1 port map( A => n12, Z => net56070);
   U85 : BUF_X1 port map( A => n7, Z => net56040);
   U86 : BUF_X1 port map( A => n13, Z => net56072);
   U87 : BUF_X1 port map( A => n13, Z => net56074);
   U88 : BUF_X1 port map( A => n8, Z => net56044);
   U89 : BUF_X1 port map( A => n8, Z => net56042);
   U90 : BUF_X1 port map( A => n13, Z => net56076);
   U91 : BUF_X1 port map( A => n8, Z => net56046);
   U92 : AOI222_X1 port map( A1 => A(3), A2 => net56040, B1 => B(3), B2 => 
                           net56046, C1 => F(3), C2 => net56052, ZN => n31);
   U93 : AOI222_X1 port map( A1 => A(8), A2 => net56040, B1 => B(8), B2 => 
                           net56046, C1 => F(8), C2 => net56052, ZN => n16);
   U94 : AOI222_X1 port map( A1 => A(31), A2 => net56040, B1 => B(31), B2 => 
                           net56046, C1 => F(31), C2 => net56052, ZN => n34);
   U95 : AOI222_X1 port map( A1 => A(17), A2 => net56036, B1 => B(17), B2 => 
                           net56042, C1 => F(17), C2 => net56048, ZN => n82);
   U96 : AOI222_X1 port map( A1 => A(14), A2 => net56036, B1 => B(14), B2 => 
                           net56042, C1 => F(14), C2 => net56048, ZN => n91);
   U97 : AOI222_X1 port map( A1 => A(28), A2 => net56038, B1 => B(28), B2 => 
                           net56044, C1 => F(28), C2 => net56050, ZN => n46);
   U98 : AOI222_X1 port map( A1 => A(23), A2 => net56038, B1 => B(23), B2 => 
                           net56044, C1 => F(23), C2 => net56050, ZN => n61);
   U99 : AOI222_X1 port map( A1 => A(15), A2 => net56036, B1 => B(15), B2 => 
                           net56042, C1 => F(15), C2 => net56048, ZN => n88);
   U100 : AOI222_X1 port map( A1 => A(27), A2 => net56038, B1 => B(27), B2 => 
                           net56044, C1 => F(27), C2 => net56050, ZN => n49);
   U101 : AOI222_X1 port map( A1 => A(16), A2 => net56036, B1 => B(16), B2 => 
                           net56042, C1 => F(16), C2 => net56048, ZN => n85);
   U102 : AOI222_X1 port map( A1 => A(24), A2 => net56038, B1 => B(24), B2 => 
                           net56044, C1 => F(24), C2 => net56050, ZN => n58);
   U103 : AOI222_X1 port map( A1 => A(21), A2 => net56038, B1 => B(21), B2 => 
                           net56044, C1 => F(21), C2 => net56050, ZN => n67);
   U104 : AOI222_X1 port map( A1 => A(10), A2 => net56036, B1 => B(10), B2 => 
                           net56042, C1 => F(10), C2 => net56048, ZN => n103);
   U105 : AOI222_X1 port map( A1 => A(25), A2 => net56038, B1 => B(25), B2 => 
                           net56044, C1 => F(25), C2 => net56050, ZN => n55);
   U106 : AOI222_X1 port map( A1 => A(22), A2 => net56038, B1 => B(22), B2 => 
                           net56044, C1 => F(22), C2 => net56050, ZN => n64);
   U107 : AOI222_X1 port map( A1 => A(19), A2 => net56036, B1 => B(19), B2 => 
                           net56042, C1 => F(19), C2 => net56048, ZN => n76);
   U108 : AOI222_X1 port map( A1 => A(20), A2 => net56038, B1 => B(20), B2 => 
                           net56044, C1 => F(20), C2 => net56050, ZN => n70);
   U109 : AOI222_X1 port map( A1 => A(13), A2 => net56036, B1 => B(13), B2 => 
                           net56042, C1 => F(13), C2 => net56048, ZN => n94);
   U112 : AOI222_X1 port map( A1 => A(26), A2 => net56038, B1 => B(26), B2 => 
                           net56044, C1 => F(26), C2 => net56050, ZN => n52);
   U114 : AOI222_X1 port map( A1 => A(29), A2 => net56038, B1 => B(29), B2 => 
                           net56044, C1 => F(29), C2 => net56050, ZN => n43);
   U117 : AOI222_X1 port map( A1 => A(30), A2 => net56038, B1 => B(30), B2 => 
                           net56044, C1 => F(30), C2 => net56050, ZN => n37);
   U138 : AOI22_X1 port map( A1 => D(5), A2 => net56058, B1 => H(5), B2 => 
                           net56064, ZN => n24);
   U139 : AOI22_X1 port map( A1 => E(0), A2 => net56066, B1 => C(0), B2 => 
                           net56072, ZN => n104);
   U141 : AOI22_X1 port map( A1 => D(31), A2 => net56058, B1 => H(31), B2 => 
                           net56064, ZN => n33);
   U142 : AOI22_X1 port map( A1 => D(12), A2 => net56054, B1 => H(12), B2 => 
                           net56060, ZN => n96);
   U143 : AOI22_X1 port map( A1 => D(28), A2 => net56056, B1 => H(28), B2 => 
                           net56062, ZN => n45);
   U144 : AOI22_X1 port map( A1 => D(30), A2 => net56056, B1 => H(30), B2 => 
                           net56062, ZN => n36);
   U145 : AOI22_X1 port map( A1 => D(7), A2 => net56058, B1 => H(7), B2 => 
                           net56064, ZN => n18);
   U146 : AOI22_X1 port map( A1 => D(17), A2 => net56054, B1 => H(17), B2 => 
                           net56060, ZN => n81);
   U147 : AOI22_X1 port map( A1 => D(2), A2 => net56056, B1 => H(2), B2 => 
                           net56062, ZN => n39);
   U148 : AOI22_X1 port map( A1 => D(21), A2 => net56056, B1 => H(21), B2 => 
                           net56062, ZN => n66);
   U149 : AOI22_X1 port map( A1 => D(9), A2 => net56058, B1 => H(9), B2 => 
                           net56064, ZN => n5);
   U150 : AOI22_X1 port map( A1 => D(14), A2 => net56054, B1 => H(14), B2 => 
                           net56060, ZN => n90);
   U151 : AOI22_X1 port map( A1 => D(6), A2 => net56058, B1 => H(6), B2 => 
                           net56064, ZN => n21);
   U152 : AOI22_X1 port map( A1 => D(20), A2 => net56056, B1 => H(20), B2 => 
                           net56062, ZN => n69);
   U153 : AOI22_X1 port map( A1 => D(4), A2 => net56058, B1 => H(4), B2 => 
                           net56064, ZN => n27);
   U154 : AOI22_X1 port map( A1 => D(23), A2 => net56056, B1 => H(23), B2 => 
                           net56062, ZN => n60);
   U155 : AOI22_X1 port map( A1 => D(11), A2 => net56054, B1 => H(11), B2 => 
                           net56060, ZN => n99);
   U156 : AOI22_X1 port map( A1 => D(18), A2 => net56054, B1 => H(18), B2 => 
                           net56060, ZN => n78);
   U157 : AOI22_X1 port map( A1 => D(29), A2 => net56056, B1 => H(29), B2 => 
                           net56062, ZN => n42);
   U158 : AOI22_X1 port map( A1 => D(1), A2 => net56054, B1 => H(1), B2 => 
                           net56060, ZN => n72);
   U159 : AOI22_X1 port map( A1 => D(15), A2 => net56054, B1 => H(15), B2 => 
                           net56060, ZN => n87);
   U160 : AOI22_X1 port map( A1 => D(25), A2 => net56056, B1 => H(25), B2 => 
                           net56062, ZN => n54);
   U161 : AOI22_X1 port map( A1 => D(27), A2 => net56056, B1 => H(27), B2 => 
                           net56062, ZN => n48);
   U162 : AOI22_X1 port map( A1 => D(26), A2 => net56056, B1 => H(26), B2 => 
                           net56062, ZN => n51);
   U163 : AOI22_X1 port map( A1 => D(16), A2 => net56054, B1 => H(16), B2 => 
                           net56060, ZN => n84);
   U164 : AOI22_X1 port map( A1 => D(24), A2 => net56056, B1 => H(24), B2 => 
                           net56062, ZN => n57);
   U165 : AOI22_X1 port map( A1 => D(10), A2 => net56054, B1 => H(10), B2 => 
                           net56060, ZN => n102);
   U166 : AOI22_X1 port map( A1 => D(3), A2 => net56058, B1 => H(3), B2 => 
                           net56064, ZN => n30);
   U167 : AOI22_X1 port map( A1 => D(22), A2 => net56056, B1 => H(22), B2 => 
                           net56062, ZN => n63);
   U168 : AOI22_X1 port map( A1 => D(19), A2 => net56054, B1 => H(19), B2 => 
                           net56060, ZN => n75);
   U169 : AOI22_X1 port map( A1 => D(8), A2 => net56058, B1 => H(8), B2 => 
                           net56064, ZN => n15);
   U170 : AOI22_X1 port map( A1 => D(13), A2 => net56054, B1 => H(13), B2 => 
                           net56060, ZN => n93);
   U171 : AOI22_X1 port map( A1 => E(6), A2 => net56070, B1 => C(6), B2 => 
                           net56076, ZN => n20);
   U172 : AOI22_X1 port map( A1 => E(7), A2 => net56070, B1 => C(7), B2 => 
                           net56076, ZN => n17);
   U173 : AOI22_X1 port map( A1 => E(9), A2 => net56070, B1 => C(9), B2 => 
                           net56076, ZN => n4);
   U174 : AOI22_X1 port map( A1 => E(8), A2 => net56070, B1 => C(8), B2 => 
                           net56076, ZN => n14);
   U175 : AOI22_X1 port map( A1 => E(5), A2 => net56070, B1 => C(5), B2 => 
                           net56076, ZN => n23);
   U176 : AOI22_X1 port map( A1 => E(3), A2 => net56070, B1 => C(3), B2 => 
                           net56076, ZN => n29);
   U177 : AOI22_X1 port map( A1 => E(30), A2 => net56068, B1 => C(30), B2 => 
                           net56074, ZN => n35);
   U178 : AOI22_X1 port map( A1 => E(21), A2 => net56068, B1 => C(21), B2 => 
                           net56074, ZN => n65);
   U179 : AOI22_X1 port map( A1 => E(28), A2 => net56068, B1 => C(28), B2 => 
                           net56074, ZN => n44);
   U180 : AOI22_X1 port map( A1 => E(20), A2 => net56068, B1 => C(20), B2 => 
                           net56074, ZN => n68);
   U181 : AOI22_X1 port map( A1 => E(29), A2 => net56068, B1 => C(29), B2 => 
                           net56074, ZN => n41);
   U182 : AOI22_X1 port map( A1 => E(25), A2 => net56068, B1 => C(25), B2 => 
                           net56074, ZN => n53);
   U183 : AOI22_X1 port map( A1 => E(26), A2 => net56068, B1 => C(26), B2 => 
                           net56074, ZN => n50);
   U184 : AOI22_X1 port map( A1 => E(27), A2 => net56068, B1 => C(27), B2 => 
                           net56074, ZN => n47);
   U185 : AOI22_X1 port map( A1 => E(22), A2 => net56068, B1 => C(22), B2 => 
                           net56074, ZN => n62);
   U186 : AOI22_X1 port map( A1 => E(2), A2 => net56068, B1 => C(2), B2 => 
                           net56074, ZN => n38);
   U187 : AOI22_X1 port map( A1 => E(23), A2 => net56068, B1 => C(23), B2 => 
                           net56074, ZN => n59);
   U188 : AOI22_X1 port map( A1 => E(24), A2 => net56068, B1 => C(24), B2 => 
                           net56074, ZN => n56);
   U189 : AOI22_X1 port map( A1 => E(15), A2 => net56066, B1 => C(15), B2 => 
                           net56072, ZN => n86);
   U190 : AOI22_X1 port map( A1 => E(10), A2 => net56066, B1 => C(10), B2 => 
                           net56072, ZN => n101);
   U191 : AOI22_X1 port map( A1 => E(13), A2 => net56066, B1 => C(13), B2 => 
                           net56072, ZN => n92);
   U192 : AOI22_X1 port map( A1 => E(14), A2 => net56066, B1 => C(14), B2 => 
                           net56072, ZN => n89);
   U193 : AOI22_X1 port map( A1 => E(11), A2 => net56066, B1 => C(11), B2 => 
                           net56072, ZN => n98);
   U194 : AOI22_X1 port map( A1 => E(16), A2 => net56066, B1 => C(16), B2 => 
                           net56072, ZN => n83);
   U195 : AOI22_X1 port map( A1 => E(12), A2 => net56066, B1 => C(12), B2 => 
                           net56072, ZN => n95);
   U196 : AOI22_X1 port map( A1 => E(17), A2 => net56066, B1 => C(17), B2 => 
                           net56072, ZN => n80);
   U197 : AOI22_X1 port map( A1 => E(18), A2 => net56066, B1 => C(18), B2 => 
                           net56072, ZN => n77);
   U198 : AOI22_X1 port map( A1 => E(19), A2 => net56066, B1 => C(19), B2 => 
                           net56072, ZN => n74);
   U199 : AOI22_X1 port map( A1 => E(1), A2 => net56066, B1 => C(1), B2 => 
                           net56072, ZN => n71);
   U200 : NOR2_X1 port map( A1 => sel(2), A2 => sel(3), ZN => n108);
   U201 : NOR2_X1 port map( A1 => n153, A2 => sel(3), ZN => n107);
   U202 : INV_X1 port map( A => sel(2), ZN => n153);
   U203 : INV_X1 port map( A => sel(0), ZN => net52587);
   U204 : AOI22_X1 port map( A1 => E(31), A2 => net56070, B1 => C(31), B2 => 
                           net56076, ZN => n32);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity comparator is

   port( r1, r2 : in std_logic_vector (31 downto 0);  sel : in std_logic_vector
         (2 downto 0);  data_out : out std_logic_vector (31 downto 0));

end comparator;

architecture SYN_beh of comparator is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, N26, N27, N28, data_out_0_port, n1, n5, n6, n8, 
      net52585, n7, n9, n10, n11, n12, n13, n_1124, n_1125, n_1126 : std_logic;

begin
   data_out <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      data_out_0_port );
   
   X_Logic0_port <= '0';
   n1 <= '0';
   r69 : comparator_DW01_cmp6_0 port map( A(31) => r1(31), A(30) => r1(30), 
                           A(29) => r1(29), A(28) => r1(28), A(27) => r1(27), 
                           A(26) => r1(26), A(25) => r1(25), A(24) => r1(24), 
                           A(23) => r1(23), A(22) => r1(22), A(21) => r1(21), 
                           A(20) => r1(20), A(19) => r1(19), A(18) => r1(18), 
                           A(17) => r1(17), A(16) => r1(16), A(15) => r1(15), 
                           A(14) => r1(14), A(13) => r1(13), A(12) => r1(12), 
                           A(11) => r1(11), A(10) => r1(10), A(9) => r1(9), 
                           A(8) => r1(8), A(7) => r1(7), A(6) => r1(6), A(5) =>
                           r1(5), A(4) => r1(4), A(3) => r1(3), A(2) => r1(2), 
                           A(1) => r1(1), A(0) => r1(0), B(31) => r2(31), B(30)
                           => r2(30), B(29) => r2(29), B(28) => r2(28), B(27) 
                           => r2(27), B(26) => r2(26), B(25) => r2(25), B(24) 
                           => r2(24), B(23) => r2(23), B(22) => r2(22), B(21) 
                           => r2(21), B(20) => r2(20), B(19) => r2(19), B(18) 
                           => r2(18), B(17) => r2(17), B(16) => r2(16), B(15) 
                           => r2(15), B(14) => r2(14), B(13) => r2(13), B(12) 
                           => r2(12), B(11) => r2(11), B(10) => r2(10), B(9) =>
                           r2(9), B(8) => r2(8), B(7) => r2(7), B(6) => r2(6), 
                           B(5) => r2(5), B(4) => r2(4), B(3) => r2(3), B(2) =>
                           r2(2), B(1) => r2(1), B(0) => r2(0), TC => n1, LT =>
                           n_1124, GT => n_1125, EQ => N26, LE => N27, GE => 
                           N28, NE => n_1126);
   U2 : NAND2_X1 port map( A1 => N26, A2 => n7, ZN => n9);
   U4 : NAND2_X1 port map( A1 => N27, A2 => sel(0), ZN => n10);
   U5 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => net52585);
   U6 : INV_X1 port map( A => sel(0), ZN => n7);
   U7 : OR2_X1 port map( A1 => n12, A2 => n11, ZN => n6);
   U8 : NAND2_X1 port map( A1 => sel(2), A2 => n13, ZN => n11);
   U9 : XNOR2_X1 port map( A => N28, B => n7, ZN => n8);
   U10 : MUX2_X1 port map( A => N27, B => N26, S => n7, Z => n12);
   U11 : AOI22_X1 port map( A1 => sel(1), A2 => n8, B1 => net52585, B2 => n13, 
                           ZN => n5);
   U12 : INV_X1 port map( A => sel(1), ZN => n13);
   U13 : OAI21_X1 port map( B1 => n5, B2 => sel(2), A => n6, ZN => 
                           data_out_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity shifter_dx_nbit32 is

   port( r1, r2 : in std_logic_vector (31 downto 0);  log : in std_logic;  
         data_out : out std_logic_vector (31 downto 0));

end shifter_dx_nbit32;

architecture SYN_beh of shifter_dx_nbit32 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069,
      N2070, N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079, 
      N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089, 
      N2090, N2091, n1, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
      n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, 
      n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
      n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
      n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, 
      n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, 
      n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803 : std_logic;

begin
   
   data_out_reg_31_inst : DLH_X1 port map( G => n1, D => N2091, Q => 
                           data_out(31));
   data_out_reg_30_inst : DLH_X1 port map( G => n1, D => N2090, Q => 
                           data_out(30));
   data_out_reg_29_inst : DLH_X1 port map( G => n1, D => N2089, Q => 
                           data_out(29));
   data_out_reg_28_inst : DLH_X1 port map( G => n1, D => N2088, Q => 
                           data_out(28));
   data_out_reg_27_inst : DLH_X1 port map( G => n1, D => N2087, Q => 
                           data_out(27));
   data_out_reg_26_inst : DLH_X1 port map( G => n1, D => N2086, Q => 
                           data_out(26));
   data_out_reg_25_inst : DLH_X1 port map( G => n1, D => N2085, Q => 
                           data_out(25));
   data_out_reg_24_inst : DLH_X1 port map( G => n1, D => N2084, Q => 
                           data_out(24));
   data_out_reg_23_inst : DLH_X1 port map( G => n1, D => N2083, Q => 
                           data_out(23));
   data_out_reg_22_inst : DLH_X1 port map( G => n1, D => N2082, Q => 
                           data_out(22));
   data_out_reg_21_inst : DLH_X1 port map( G => n1, D => N2081, Q => 
                           data_out(21));
   data_out_reg_20_inst : DLH_X1 port map( G => n1, D => N2080, Q => 
                           data_out(20));
   data_out_reg_19_inst : DLH_X1 port map( G => n1, D => N2079, Q => 
                           data_out(19));
   data_out_reg_18_inst : DLH_X1 port map( G => n1, D => N2078, Q => 
                           data_out(18));
   data_out_reg_17_inst : DLH_X1 port map( G => n1, D => N2077, Q => 
                           data_out(17));
   data_out_reg_16_inst : DLH_X1 port map( G => n1, D => N2076, Q => 
                           data_out(16));
   data_out_reg_15_inst : DLH_X1 port map( G => n1, D => N2075, Q => 
                           data_out(15));
   data_out_reg_14_inst : DLH_X1 port map( G => n1, D => N2074, Q => 
                           data_out(14));
   data_out_reg_13_inst : DLH_X1 port map( G => n1, D => N2073, Q => 
                           data_out(13));
   data_out_reg_12_inst : DLH_X1 port map( G => n1, D => N2072, Q => 
                           data_out(12));
   data_out_reg_11_inst : DLH_X1 port map( G => n1, D => N2071, Q => 
                           data_out(11));
   data_out_reg_10_inst : DLH_X1 port map( G => n1, D => N2070, Q => 
                           data_out(10));
   data_out_reg_9_inst : DLH_X1 port map( G => n1, D => N2069, Q => data_out(9)
                           );
   data_out_reg_8_inst : DLH_X1 port map( G => n1, D => N2068, Q => data_out(8)
                           );
   data_out_reg_7_inst : DLH_X1 port map( G => n1, D => N2067, Q => data_out(7)
                           );
   data_out_reg_6_inst : DLH_X1 port map( G => n1, D => N2066, Q => data_out(6)
                           );
   data_out_reg_5_inst : DLH_X1 port map( G => n1, D => N2065, Q => data_out(5)
                           );
   data_out_reg_4_inst : DLH_X1 port map( G => n1, D => N2064, Q => data_out(4)
                           );
   data_out_reg_3_inst : DLH_X1 port map( G => n1, D => N2063, Q => data_out(3)
                           );
   data_out_reg_2_inst : DLH_X1 port map( G => n1, D => N2062, Q => data_out(2)
                           );
   data_out_reg_1_inst : DLH_X1 port map( G => n1, D => N2061, Q => data_out(1)
                           );
   data_out_reg_0_inst : DLH_X1 port map( G => n1, D => N2060, Q => data_out(0)
                           );
   n1 <= '1';
   U367 : NAND2_X2 port map( A1 => n481, A2 => n489, ZN => n284);
   U392 : NAND2_X2 port map( A1 => n482, A2 => n652, ZN => n196);
   U408 : AND3_X2 port map( A1 => n774, A2 => n798, A3 => r2(4), ZN => n479);
   U524 : NAND3_X1 port map( A1 => n123, A2 => n124, A3 => n125, ZN => n121);
   U525 : NAND3_X1 port map( A1 => n746, A2 => n135, A3 => n626, ZN => n131);
   U526 : NAND3_X1 port map( A1 => n659, A2 => n661, A3 => n140, ZN => n139);
   U527 : NAND3_X1 port map( A1 => n656, A2 => n662, A3 => r1(25), ZN => n156);
   U528 : NAND3_X1 port map( A1 => n179, A2 => n180, A3 => n181, ZN => N2080);
   U529 : NAND3_X1 port map( A1 => n761, A2 => n185, A3 => n186, ZN => n184);
   U530 : NAND3_X1 port map( A1 => n187, A2 => n188, A3 => n189, ZN => n182);
   U531 : NAND3_X1 port map( A1 => n203, A2 => n204, A3 => n205, ZN => n199);
   U533 : NAND3_X1 port map( A1 => n314, A2 => n315, A3 => n316, ZN => N2070);
   U534 : NAND3_X1 port map( A1 => n373, A2 => n374, A3 => n375, ZN => n369);
   U535 : NAND3_X1 port map( A1 => n419, A2 => n420, A3 => n421, ZN => N2063);
   U536 : NAND3_X1 port map( A1 => n425, A2 => n427, A3 => n426, ZN => n424);
   U537 : NAND3_X1 port map( A1 => n435, A2 => n436, A3 => n437, ZN => N2062);
   U538 : NAND3_X1 port map( A1 => n763, A2 => n105, A3 => log, ZN => n158);
   U539 : NAND3_X1 port map( A1 => n450, A2 => n751, A3 => n451, ZN => N2061);
   U540 : NAND3_X1 port map( A1 => n372, A2 => n387, A3 => n371, ZN => n334);
   U3 : INV_X1 port map( A => n780, ZN => n553);
   U4 : INV_X2 port map( A => n227, ZN => n781);
   U5 : AND3_X2 port map( A1 => r2(0), A2 => n774, A3 => r2(4), ZN => n481);
   U6 : OAI222_X1 port map( A1 => n695, A2 => n646, B1 => n697, B2 => n644, C1 
                           => n656, C2 => n801, ZN => n292);
   U7 : OAI221_X1 port map( B1 => n654, B2 => n665, C1 => n196, C2 => n676, A 
                           => n467, ZN => n463);
   U8 : OAI222_X1 port map( A1 => n646, A2 => n691, B1 => n695, B2 => n644, C1 
                           => n655, C2 => n679, ZN => n310);
   U9 : NOR3_X1 port map( A1 => n796, A2 => r2(1), A3 => n795, ZN => n482);
   U10 : BUF_X1 port map( A => n498, Z => n652);
   U11 : NOR3_X1 port map( A1 => r2(1), A2 => r2(2), A3 => n795, ZN => n483);
   U12 : BUF_X1 port map( A => n608, Z => n653);
   U13 : INV_X1 port map( A => n624, ZN => n230);
   U14 : NAND2_X1 port map( A1 => n482, A2 => n606, ZN => n227);
   U15 : OAI222_X1 port map( A1 => n699, A2 => n285, B1 => n412, B2 => n605, C1
                           => n697, C2 => n284, ZN => n410);
   U16 : OR2_X1 port map( A1 => n297, A2 => n775, ZN => n620);
   U17 : AND2_X1 port map( A1 => n575, A2 => n576, ZN => n174);
   U18 : INV_X1 port map( A => n566, ZN => n106);
   U19 : OR2_X2 port map( A1 => n582, A2 => n334, ZN => n566);
   U20 : INV_X1 port map( A => n571, ZN => n98);
   U21 : BUF_X1 port map( A => n176, Z => n607);
   U22 : AND3_X1 port map( A1 => n397, A2 => n396, A3 => n395, ZN => n554);
   U23 : OR3_X1 port map( A1 => n361, A2 => n363, A3 => n362, ZN => n555);
   U24 : OR3_X1 port map( A1 => n310, A2 => n312, A3 => n311, ZN => n556);
   U25 : OR3_X1 port map( A1 => n465, A2 => n464, A3 => n466, ZN => n557);
   U26 : OR3_X1 port map( A1 => n292, A2 => n293, A3 => n294, ZN => n558);
   U27 : OR3_X1 port map( A1 => n415, A2 => n416, A3 => n414, ZN => n559);
   U28 : AND2_X1 port map( A1 => n304, A2 => n301, ZN => n560);
   U29 : OR3_X1 port map( A1 => r2(17), A2 => r2(18), A3 => r2(16), ZN => n561)
                           ;
   U30 : OR3_X1 port map( A1 => r2(24), A2 => r2(25), A3 => r2(23), ZN => n562)
                           ;
   U31 : OR2_X1 port map( A1 => n798, A2 => r2(4), ZN => n563);
   U32 : AND2_X1 port map( A1 => n594, A2 => n593, ZN => n564);
   U33 : OR2_X1 port map( A1 => n753, A2 => n756, ZN => n565);
   U34 : NOR2_X1 port map( A1 => n281, A2 => n565, ZN => n280);
   U35 : BUF_X2 port map( A => n168, Z => n646);
   U36 : BUF_X2 port map( A => n197, Z => n644);
   U37 : AOI221_X1 port map( B1 => r1(20), B2 => n788, C1 => r1(19), C2 => n107
                           , A => n791, ZN => n236);
   U38 : NOR2_X1 port map( A1 => n413, A2 => n559, ZN => n412);
   U39 : NOR3_X1 port map( A1 => n567, A2 => n568, A3 => n569, ZN => n441);
   U40 : NAND3_X1 port map( A1 => n622, A2 => n621, A3 => n623, ZN => n567);
   U41 : AND2_X1 port map( A1 => n760, A2 => n683, ZN => n568);
   U42 : AND2_X1 port map( A1 => n790, A2 => n680, ZN => n569);
   U43 : CLKBUF_X1 port map( A => n763, Z => n570);
   U44 : NAND2_X1 port map( A1 => n479, A2 => n489, ZN => n270);
   U45 : NAND2_X1 port map( A1 => n479, A2 => n497, ZN => n285);
   U46 : NAND2_X2 port map( A1 => n479, A2 => n491, ZN => n249);
   U47 : AND2_X1 port map( A1 => n491, A2 => n653, ZN => n571);
   U48 : BUF_X1 port map( A => n490, Z => n606);
   U49 : AND3_X2 port map( A1 => n477, A2 => n476, A3 => n407, ZN => n371);
   U50 : NAND3_X1 port map( A1 => n207, A2 => n215, A3 => n107, ZN => n572);
   U51 : NAND3_X1 port map( A1 => n207, A2 => n215, A3 => n107, ZN => n573);
   U52 : INV_X1 port map( A => n145, ZN => n574);
   U53 : AND2_X1 port map( A1 => n499, A2 => n652, ZN => n625);
   U54 : BUF_X1 port map( A => n490, Z => n650);
   U55 : NOR2_X1 port map( A1 => n647, A2 => n563, ZN => n490);
   U56 : NAND2_X1 port map( A1 => n185, A2 => n186, ZN => n575);
   U57 : INV_X1 port map( A => n157, ZN => n576);
   U58 : INV_X1 port map( A => n582, ZN => n185);
   U59 : NAND2_X1 port map( A1 => n398, A2 => n554, ZN => n394);
   U60 : AOI221_X1 port map( B1 => n688, B2 => n788, C1 => r1(20), C2 => n107, 
                           A => n791, ZN => n221);
   U61 : NAND2_X1 port map( A1 => n306, A2 => n560, ZN => n299);
   U62 : OR2_X1 port map( A1 => n98, A2 => n673, ZN => n577);
   U63 : OR2_X1 port map( A1 => n101, A2 => n803, ZN => n578);
   U64 : NAND3_X1 port map( A1 => n577, A2 => n578, A3 => n298, ZN => N2071);
   U65 : BUF_X1 port map( A => n127, Z => n579);
   U66 : AND2_X1 port map( A1 => n715, A2 => n600, ZN => n580);
   U67 : AND2_X1 port map( A1 => n725, A2 => n601, ZN => n581);
   U68 : NOR3_X1 port map( A1 => n580, A2 => n581, A3 => n749, ZN => n110);
   U69 : NAND2_X1 port map( A1 => n278, A2 => n564, ZN => N2072);
   U70 : OR3_X2 port map( A1 => n755, A2 => n767, A3 => n296, ZN => n582);
   U71 : AOI21_X2 port map( B1 => n582, B2 => n736, A => n264, ZN => n163);
   U72 : AND2_X1 port map( A1 => n680, A2 => n600, ZN => n583);
   U73 : AND2_X1 port map( A1 => n624, A2 => n776, ZN => n584);
   U74 : NOR3_X1 port map( A1 => n225, A2 => n584, A3 => n583, ZN => n224);
   U75 : CLKBUF_X3 port map( A => n572, Z => n654);
   U76 : BUF_X1 port map( A => n145, Z => n649);
   U77 : OAI221_X1 port map( B1 => n654, B2 => n668, C1 => n196, C2 => n800, A 
                           => n417, ZN => n413);
   U78 : NAND2_X1 port map( A1 => n369, A2 => n268, ZN => n585);
   U79 : NAND2_X1 port map( A1 => n737, A2 => n370, ZN => n586);
   U80 : AND3_X1 port map( A1 => n585, A2 => n586, A3 => n751, ZN => n368);
   U81 : NAND2_X1 port map( A1 => n770, A2 => n700, ZN => n587);
   U82 : NAND2_X1 port map( A1 => n214, A2 => n377, ZN => n588);
   U83 : NAND2_X1 port map( A1 => n759, A2 => n704, ZN => n589);
   U84 : AND3_X1 port map( A1 => n587, A2 => n588, A3 => n589, ZN => n374);
   U85 : BUF_X2 port map( A => n490, Z => n651);
   U86 : NOR2_X1 port map( A1 => n463, A2 => n557, ZN => n462);
   U87 : OR2_X1 port map( A1 => n691, A2 => n285, ZN => n590);
   U88 : OR2_X1 port map( A1 => n462, A2 => n605, ZN => n591);
   U89 : OR2_X1 port map( A1 => n802, A2 => n284, ZN => n592);
   U90 : NAND3_X1 port map( A1 => n590, A2 => n591, A3 => n592, ZN => n460);
   U91 : OR2_X1 port map( A1 => n98, A2 => n803, ZN => n593);
   U92 : OR2_X1 port map( A1 => n101, A2 => n676, ZN => n594);
   U93 : INV_X1 port map( A => n601, ZN => n101);
   U94 : NOR2_X1 port map( A1 => n360, A2 => n555, ZN => n359);
   U95 : AND2_X1 port map( A1 => n790, A2 => n694, ZN => n595);
   U96 : AND2_X1 port map( A1 => n760, A2 => n696, ZN => n596);
   U97 : NOR3_X1 port map( A1 => n595, A2 => n596, A3 => n358, ZN => n357);
   U98 : OAI222_X1 port map( A1 => n802, A2 => n285, B1 => n487, B2 => n605, C1
                           => n799, C2 => n284, ZN => n485);
   U99 : OAI221_X1 port map( B1 => n654, B2 => n664, C1 => n196, C2 => n803, A 
                           => n496, ZN => n492);
   U100 : NOR2_X1 port map( A1 => n309, A2 => n556, ZN => n308);
   U101 : OR2_X1 port map( A1 => n707, A2 => n247, ZN => n597);
   U102 : OR2_X1 port map( A1 => n308, A2 => n222, ZN => n598);
   U103 : OR2_X1 port map( A1 => n712, A2 => n249, ZN => n599);
   U104 : NAND3_X1 port map( A1 => n597, A2 => n598, A3 => n599, ZN => n305);
   U105 : NAND2_X1 port map( A1 => n249, A2 => n247, ZN => n222);
   U106 : AND2_X1 port map( A1 => n284, A2 => n285, ZN => n488);
   U107 : INV_X1 port map( A => n284, ZN => n770);
   U108 : INV_X1 port map( A => n285, ZN => n759);
   U109 : BUF_X1 port map( A => n641, Z => n642);
   U110 : INV_X2 port map( A => n98, ZN => n600);
   U111 : AND2_X4 port map( A1 => n651, A2 => n491, ZN => n601);
   U112 : OR4_X2 port map( A1 => r2(7), A2 => r2(6), A3 => r2(8), A4 => r2(9), 
                           ZN => n505);
   U113 : OR4_X1 port map( A1 => r2(27), A2 => r2(26), A3 => r2(29), A4 => 
                           r2(28), ZN => n506);
   U114 : NOR2_X1 port map( A1 => n507, A2 => n561, ZN => n502);
   U115 : NOR2_X1 port map( A1 => n291, A2 => n558, ZN => n290);
   U116 : OR2_X1 port map( A1 => n712, A2 => n247, ZN => n602);
   U117 : OR2_X1 port map( A1 => n290, A2 => n222, ZN => n603);
   U118 : OR2_X1 port map( A1 => n718, A2 => n249, ZN => n604);
   U119 : NAND3_X1 port map( A1 => n602, A2 => n603, A3 => n604, ZN => n288);
   U120 : OR4_X1 port map( A1 => r2(20), A2 => r2(19), A3 => r2(22), A4 => 
                           r2(21), ZN => n507);
   U121 : NAND2_X2 port map( A1 => n480, A2 => n651, ZN => n247);
   U122 : INV_X1 port map( A => n625, ZN => n145);
   U123 : OR2_X2 port map( A1 => n222, A2 => n582, ZN => n605);
   U124 : NOR3_X1 port map( A1 => r2(0), A2 => r2(4), A3 => n647, ZN => n608);
   U125 : NOR3_X1 port map( A1 => r2(0), A2 => r2(4), A3 => n647, ZN => n498);
   U126 : INV_X2 port map( A => n793, ZN => n640);
   U127 : INV_X1 port map( A => n227, ZN => n609);
   U128 : NAND2_X1 port map( A1 => n608, A2 => n483, ZN => n177);
   U129 : OR2_X1 port map( A1 => n713, A2 => n285, ZN => n610);
   U130 : OR2_X1 port map( A1 => n359, A2 => n605, ZN => n611);
   U131 : OR2_X1 port map( A1 => n706, A2 => n284, ZN => n612);
   U132 : NAND3_X1 port map( A1 => n610, A2 => n611, A3 => n612, ZN => n358);
   U133 : OAI221_X1 port map( B1 => n654, B2 => n671, C1 => n196, C2 => n799, A
                           => n364, ZN => n360);
   U134 : OR2_X1 port map( A1 => n98, A2 => n667, ZN => n613);
   U135 : OR2_X1 port map( A1 => n101, A2 => n668, ZN => n614);
   U136 : NAND3_X1 port map( A1 => n613, A2 => n614, A3 => n383, ZN => N2065);
   U137 : NAND2_X1 port map( A1 => n123, A2 => n384, ZN => n615);
   U138 : NAND2_X1 port map( A1 => n385, A2 => n776, ZN => n616);
   U139 : AND3_X1 port map( A1 => n615, A2 => n616, A3 => n751, ZN => n383);
   U140 : NOR3_X1 port map( A1 => n601, A2 => n571, A3 => n648, ZN => n123);
   U141 : AND2_X1 port map( A1 => r1(9), A2 => n600, ZN => n617);
   U142 : AND2_X1 port map( A1 => n333, A2 => n745, ZN => n618);
   U143 : AND2_X1 port map( A1 => n758, A2 => n776, ZN => n619);
   U144 : NOR3_X1 port map( A1 => n617, A2 => n618, A3 => n619, ZN => n328);
   U145 : NAND2_X1 port map( A1 => n105, A2 => n752, ZN => n297);
   U146 : OR2_X1 port map( A1 => n695, A2 => n285, ZN => n621);
   U147 : OR2_X1 port map( A1 => n443, A2 => n605, ZN => n622);
   U148 : OR2_X1 port map( A1 => n691, A2 => n284, ZN => n623);
   U149 : OAI221_X1 port map( B1 => n654, B2 => n666, C1 => n196, C2 => n679, A
                           => n448, ZN => n444);
   U150 : AND2_X4 port map( A1 => n480, A2 => n653, ZN => n624);
   U151 : BUF_X1 port map( A => n99, Z => n648);
   U152 : BUF_X1 port map( A => n153, Z => n641);
   U153 : AND3_X1 port map( A1 => n643, A2 => n645, A3 => n196, ZN => n207);
   U154 : INV_X1 port map( A => n643, ZN => n779);
   U155 : INV_X1 port map( A => n645, ZN => n791);
   U156 : NOR3_X1 port map( A1 => r2(1), A2 => r2(3), A3 => n796, ZN => n497);
   U157 : NOR3_X1 port map( A1 => r2(2), A2 => r2(3), A3 => n797, ZN => n489);
   U158 : NOR3_X1 port map( A1 => r2(2), A2 => r2(3), A3 => r2(1), ZN => n491);
   U159 : NOR3_X1 port map( A1 => n796, A2 => r2(3), A3 => n797, ZN => n499);
   U160 : NAND2_X1 port map( A1 => n650, A2 => n483, ZN => n176);
   U161 : NOR3_X1 port map( A1 => n786, A2 => n574, A3 => n150, ZN => n626);
   U162 : OR2_X1 port map( A1 => n733, A2 => n372, ZN => n627);
   U163 : OR2_X1 port map( A1 => n722, A2 => n387, ZN => n628);
   U164 : NAND3_X1 port map( A1 => n627, A2 => n628, A3 => n388, ZN => n384);
   U165 : NAND2_X1 port map( A1 => r1(7), A2 => n600, ZN => n629);
   U166 : NAND2_X1 port map( A1 => n762, A2 => n736, ZN => n630);
   U167 : INV_X1 port map( A => n355, ZN => n631);
   U168 : AND3_X1 port map( A1 => n629, A2 => n630, A3 => n631, ZN => n354);
   U169 : OR2_X1 port map( A1 => n802, A2 => n247, ZN => n632);
   U170 : OR2_X1 port map( A1 => n691, A2 => n249, ZN => n633);
   U171 : NAND3_X1 port map( A1 => n632, A2 => n633, A3 => n393, ZN => n389);
   U172 : NAND2_X1 port map( A1 => r1(7), A2 => n778, ZN => n634);
   U173 : NAND2_X1 port map( A1 => n680, A2 => n792, ZN => n635);
   U174 : INV_X1 port map( A => n399, ZN => n636);
   U175 : AND3_X1 port map( A1 => n634, A2 => n635, A3 => n636, ZN => n398);
   U176 : INV_X1 port map( A => n196, ZN => n792);
   U177 : NOR2_X1 port map( A1 => n506, A2 => n562, ZN => n503);
   U178 : NAND2_X1 port map( A1 => n770, A2 => n698, ZN => n637);
   U179 : NAND2_X1 port map( A1 => n214, A2 => n394, ZN => n638);
   U180 : NAND2_X1 port map( A1 => n759, A2 => n700, ZN => n639);
   U181 : AND3_X1 port map( A1 => n637, A2 => n638, A3 => n639, ZN => n393);
   U182 : NOR2_X1 port map( A1 => n105, A2 => n100, ZN => n162);
   U183 : INV_X1 port map( A => r1(24), ZN => n699);
   U184 : INV_X1 port map( A => n119, ZN => n761);
   U185 : INV_X1 port map( A => n215, ZN => n780);
   U186 : NOR2_X1 port map( A1 => n781, A2 => n624, ZN => n215);
   U187 : NAND2_X1 port map( A1 => n202, A2 => n207, ZN => n119);
   U188 : INV_X1 port map( A => n116, ZN => n742);
   U189 : INV_X1 port map( A => n282, ZN => n756);
   U190 : NOR3_X1 port map( A1 => n769, A2 => n768, A3 => n758, ZN => n282);
   U191 : NOR2_X1 port map( A1 => n222, A2 => n582, ZN => n214);
   U192 : NOR2_X1 port map( A1 => n620, A2 => n566, ZN => n157);
   U193 : OAI21_X1 port map( B1 => n163, B2 => n620, A => n751, ZN => n116);
   U194 : INV_X1 port map( A => n318, ZN => n776);
   U195 : INV_X1 port map( A => n607, ZN => n787);
   U196 : NOR2_X1 port map( A1 => n780, A2 => n222, ZN => n202);
   U197 : OAI21_X1 port map( B1 => n620, B2 => n404, A => n751, ZN => n423);
   U198 : INV_X1 port map( A => n247, ZN => n790);
   U199 : INV_X1 port map( A => n334, ZN => n763);
   U200 : INV_X1 port map( A => n123, ZN => n775);
   U201 : INV_X1 port map( A => n343, ZN => n748);
   U202 : INV_X1 port map( A => n268, ZN => n747);
   U203 : INV_X1 port map( A => n454, ZN => n766);
   U204 : INV_X1 port map( A => n730, ZN => n733);
   U205 : INV_X1 port map( A => n138, ZN => n794);
   U206 : INV_X1 port map( A => n137, ZN => n789);
   U207 : INV_X1 port map( A => n108, ZN => n788);
   U208 : AOI211_X1 port map( C1 => n761, C2 => n199, A => n201, B => n183, ZN 
                           => n200);
   U209 : OAI22_X1 port map( A1 => n722, A2 => n646, B1 => n733, B2 => n644, ZN
                           => n201);
   U210 : INV_X1 port map( A => n319, ZN => n769);
   U211 : NAND2_X1 port map( A1 => n123, A2 => n736, ZN => n318);
   U212 : INV_X1 port map( A => n332, ZN => n768);
   U213 : AOI21_X1 port map( B1 => n222, B2 => n112, A => n116, ZN => n223);
   U214 : AOI21_X1 port map( B1 => n150, B2 => n112, A => n749, ZN => n141);
   U215 : NAND4_X1 port map( A1 => n319, A2 => n332, A3 => n366, A4 => n488, ZN
                           => n296);
   U216 : AOI21_X1 port map( B1 => n296, B2 => n736, A => n264, ZN => n271);
   U217 : INV_X1 port map( A => n366, ZN => n758);
   U218 : AOI22_X1 port map( A1 => n730, A2 => n770, B1 => n737, B2 => n759, ZN
                           => n301);
   U219 : OAI21_X1 port map( B1 => n764, B2 => n772, A => n737, ZN => n404);
   U220 : NAND2_X1 port map( A1 => n123, A2 => n105, ZN => n454);
   U221 : AOI21_X1 port map( B1 => n134, B2 => n264, A => n162, ZN => n343);
   U222 : NAND2_X1 port map( A1 => n134, A2 => n570, ZN => n244);
   U223 : AOI22_X1 port map( A1 => n794, A2 => n736, B1 => n117, B2 => n118, ZN
                           => n114);
   U224 : OAI22_X1 port map( A1 => n733, A2 => n657, B1 => n784, B2 => n722, ZN
                           => n117);
   U225 : INV_X1 port map( A => n249, ZN => n760);
   U226 : INV_X1 port map( A => n387, ZN => n762);
   U227 : NAND2_X1 port map( A1 => n753, A2 => n244, ZN => n268);
   U228 : NOR3_X1 port map( A1 => n773, A2 => n764, A3 => n765, ZN => n477);
   U229 : INV_X1 port map( A => n162, ZN => n751);
   U230 : INV_X1 port map( A => n161, ZN => n749);
   U231 : AOI21_X1 port map( B1 => n127, B2 => n134, A => n162, ZN => n161);
   U232 : INV_X1 port map( A => n408, ZN => n773);
   U233 : INV_X1 port map( A => n372, ZN => n771);
   U234 : INV_X1 port map( A => n476, ZN => n772);
   U235 : CLKBUF_X1 port map( A => n108, Z => n655);
   U236 : CLKBUF_X1 port map( A => n137, Z => n658);
   U237 : CLKBUF_X1 port map( A => n138, Z => n661);
   U238 : CLKBUF_X1 port map( A => n108, Z => n656);
   U239 : CLKBUF_X1 port map( A => n137, Z => n659);
   U240 : CLKBUF_X1 port map( A => n138, Z => n662);
   U241 : CLKBUF_X1 port map( A => n108, Z => n657);
   U242 : CLKBUF_X1 port map( A => n138, Z => n663);
   U243 : CLKBUF_X1 port map( A => n137, Z => n660);
   U244 : INV_X1 port map( A => n174, ZN => n745);
   U245 : INV_X1 port map( A => n386, ZN => n765);
   U246 : NAND2_X1 port map( A1 => n229, A2 => n230, ZN => n228);
   U247 : INV_X1 port map( A => n455, ZN => n764);
   U248 : INV_X1 port map( A => n144, ZN => n746);
   U249 : INV_X1 port map( A => n118, ZN => n743);
   U250 : INV_X1 port map( A => n648, ZN => n774);
   U251 : NOR3_X1 port map( A1 => n797, A2 => n796, A3 => n795, ZN => n480);
   U252 : NOR2_X1 port map( A1 => n297, A2 => n775, ZN => n134);
   U253 : INV_X1 port map( A => n726, ZN => n722);
   U254 : NOR2_X1 port map( A1 => n576, A2 => n740, ZN => n112);
   U255 : NOR3_X1 port map( A1 => n797, A2 => r2(2), A3 => n795, ZN => n478);
   U256 : INV_X1 port map( A => n703, ZN => n700);
   U257 : AOI222_X1 port map( A1 => n768, A2 => n710, B1 => n758, B2 => n704, 
                           C1 => n769, C2 => n700, ZN => n418);
   U258 : AOI222_X1 port map( A1 => n787, A2 => n700, B1 => n779, B2 => n710, 
                           C1 => n791, C2 => n704, ZN => n240);
   U259 : INV_X1 port map( A => n690, ZN => n691);
   U260 : AOI222_X1 port map( A1 => n624, A2 => n729, B1 => n792, B2 => n715, 
                           C1 => n609, C2 => n724, ZN => n239);
   U261 : INV_X1 port map( A => n693, ZN => n695);
   U262 : NOR2_X1 port map( A1 => n738, A2 => n763, ZN => n264);
   U263 : OAI221_X1 port map( B1 => n685, B2 => n270, C1 => n682, C2 => n287, A
                           => n500, ZN => n484);
   U264 : AOI222_X1 port map( A1 => n768, A2 => n696, B1 => n758, B2 => n692, 
                           C1 => n769, C2 => n687, ZN => n500);
   U265 : AOI211_X1 port map( C1 => n783, C2 => n129, A => n566, B => n119, ZN 
                           => n126);
   U266 : INV_X1 port map( A => n124, ZN => n783);
   U267 : OAI21_X1 port map( B1 => n119, B2 => n576, A => n184, ZN => n118);
   U268 : INV_X1 port map( A => n675, ZN => n676);
   U269 : INV_X1 port map( A => n678, ZN => n679);
   U270 : AOI22_X1 port map( A1 => n761, A2 => n157, B1 => n123, B2 => n125, ZN
                           => n144);
   U271 : OAI221_X1 port map( B1 => n283, B2 => n770, C1 => n737, C2 => n284, A
                           => n285, ZN => n281);
   U272 : AOI22_X1 port map( A1 => n286, A2 => n270, B1 => n755, B2 => n733, ZN
                           => n283);
   U273 : OAI22_X1 port map( A1 => n726, A2 => n287, B1 => n288, B2 => n767, ZN
                           => n286);
   U274 : NOR3_X1 port map( A1 => n332, A2 => n738, A3 => n244, ZN => n331);
   U275 : AOI211_X1 port map( C1 => n106, C2 => n305, A => n307, B => n264, ZN 
                           => n306);
   U276 : OAI21_X1 port map( B1 => n761, B2 => n738, A => n163, ZN => n127);
   U277 : NAND2_X1 port map( A1 => n480, A2 => n481, ZN => n105);
   U278 : AOI22_X1 port map( A1 => n733, A2 => n779, B1 => n644, B2 => n198, ZN
                           => n195);
   U279 : OAI22_X1 port map( A1 => n199, A2 => n791, B1 => n646, B2 => n724, ZN
                           => n198);
   U280 : AOI22_X1 port map( A1 => r1(28), A2 => n767, B1 => n726, B2 => n755, 
                           ZN => n304);
   U281 : NAND2_X1 port map( A1 => n479, A2 => n499, ZN => n366);
   U282 : NAND2_X1 port map( A1 => n482, A2 => n479, ZN => n407);
   U283 : NAND2_X1 port map( A1 => n478, A2 => n479, ZN => n386);
   U284 : INV_X1 port map( A => r2(1), ZN => n797);
   U285 : INV_X1 port map( A => r2(2), ZN => n796);
   U286 : INV_X1 port map( A => n684, ZN => n685);
   U287 : AOI22_X1 port map( A1 => n771, A2 => n700, B1 => n762, B2 => n698, ZN
                           => n473);
   U288 : AOI22_X1 port map( A1 => n288, A2 => n106, B1 => n755, B2 => n728, ZN
                           => n289);
   U289 : AOI22_X1 port map( A1 => n789, A2 => n710, B1 => r1(26), B2 => n794, 
                           ZN => n166);
   U290 : AOI22_X1 port map( A1 => n771, A2 => n704, B1 => n762, B2 => n700, ZN
                           => n456);
   U291 : AOI22_X1 port map( A1 => n793, A2 => n710, B1 => n787, B2 => n715, ZN
                           => n204);
   U292 : AOI221_X1 port map( B1 => n696, B2 => n794, C1 => n694, C2 => n788, A
                           => n206, ZN => n205);
   U293 : OAI211_X1 port map( C1 => n740, C2 => n646, A => n169, B => n170, ZN 
                           => N2081);
   U294 : AOI22_X1 port map( A1 => n171, A2 => n761, B1 => n112, B2 => n119, ZN
                           => n169);
   U295 : AOI21_X1 port map( B1 => n172, B2 => n173, A => n174, ZN => n171);
   U296 : INV_X1 port map( A => n741, ZN => n736);
   U297 : OAI211_X1 port map( C1 => n101, C2 => n703, A => n141, B => n142, ZN 
                           => N2084);
   U298 : OAI211_X1 port map( C1 => n733, C2 => n145, A => n146, B => n147, ZN 
                           => n143);
   U299 : AOI222_X1 port map( A1 => n789, A2 => n725, B1 => r1(27), B2 => n788,
                           C1 => n794, C2 => n715, ZN => n147);
   U300 : OAI211_X1 port map( C1 => n101, C2 => n679, A => n265, B => n266, ZN 
                           => N2073);
   U301 : AOI211_X1 port map( C1 => n267, C2 => n268, A => n269, B => n162, ZN 
                           => n266);
   U302 : OAI22_X1 port map( A1 => n739, A2 => n270, B1 => n271, B2 => n620, ZN
                           => n269);
   U303 : OAI22_X1 port map( A1 => n739, A2 => n98, B1 => n648, B2 => n100, ZN 
                           => N2091);
   U304 : NAND2_X1 port map( A1 => n480, A2 => n479, ZN => n455);
   U305 : NAND2_X1 port map( A1 => n481, A2 => n483, ZN => n372);
   U306 : NOR2_X1 port map( A1 => n780, A2 => n211, ZN => n193);
   U307 : NOR2_X1 port map( A1 => n740, A2 => n282, ZN => n307);
   U308 : OAI21_X1 port map( B1 => n605, B2 => n244, A => n211, ZN => n229);
   U309 : NAND4_X1 port map( A1 => n210, A2 => n214, A3 => n553, A4 => n570, ZN
                           => n213);
   U310 : AOI21_X1 port map( B1 => n737, B2 => n406, A => n162, ZN => n405);
   U311 : OAI21_X1 port map( B1 => n297, B2 => n407, A => n408, ZN => n406);
   U312 : OAI211_X1 port map( C1 => n303, C2 => n754, A => n285, B => n284, ZN 
                           => n302);
   U313 : INV_X1 port map( A => n304, ZN => n754);
   U314 : AND3_X1 port map( A1 => n305, A2 => n287, A3 => n270, ZN => n303);
   U315 : NAND2_X1 port map( A1 => n479, A2 => n483, ZN => n387);
   U316 : AOI22_X1 port map( A1 => n793, A2 => n715, B1 => n787, B2 => n723, ZN
                           => n187);
   U317 : AOI221_X1 port map( B1 => n700, B2 => n789, C1 => n698, C2 => n794, A
                           => n190, ZN => n189);
   U318 : OAI211_X1 port map( C1 => n113, C2 => n744, A => n114, B => n115, ZN 
                           => N2087);
   U319 : INV_X1 port map( A => n112, ZN => n744);
   U320 : OAI211_X1 port map( C1 => n740, C2 => n657, A => n109, B => n110, ZN 
                           => N2088);
   U321 : NOR2_X1 port map( A1 => n743, A2 => n733, ZN => n111);
   U322 : NAND4_X1 port map( A1 => n131, A2 => n751, A3 => n132, A4 => n133, ZN
                           => N2085);
   U323 : OAI221_X1 port map( B1 => n98, B2 => n733, C1 => n740, C2 => n101, A 
                           => n102, ZN => N2090);
   U324 : BUF_X1 port map( A => n731, Z => n729);
   U325 : BUF_X1 port map( A => n732, Z => n728);
   U326 : NAND4_X1 port map( A1 => n120, A2 => n121, A3 => n751, A4 => n122, ZN
                           => N2086);
   U327 : OAI21_X1 port map( B1 => n126, B2 => n579, A => n128, ZN => n120);
   U328 : BUF_X1 port map( A => n731, Z => n730);
   U329 : INV_X1 port map( A => n186, ZN => n753);
   U330 : BUF_X1 port map( A => n732, Z => n727);
   U331 : INV_X1 port map( A => n391, ZN => n750);
   U332 : OAI222_X1 port map( A1 => n699, A2 => n247, B1 => n335, B2 => n222, 
                           C1 => n702, C2 => n249, ZN => n333);
   U333 : NOR4_X1 port map( A1 => n336, A2 => n337, A3 => n338, A4 => n339, ZN 
                           => n335);
   U334 : OAI22_X1 port map( A1 => n802, A2 => n230, B1 => n799, B2 => n227, ZN
                           => n382);
   U335 : INV_X1 port map( A => n719, ZN => n715);
   U336 : NOR4_X1 port map( A1 => n492, A2 => n493, A3 => n494, A4 => n495, ZN 
                           => n487);
   U337 : OAI222_X1 port map( A1 => n660, A2 => n667, B1 => n649, B2 => n668, 
                           C1 => n661, C2 => n666, ZN => n495);
   U338 : OAI222_X1 port map( A1 => n658, A2 => n802, B1 => n649, B2 => n691, 
                           C1 => n662, C2 => n799, ZN => n253);
   U339 : OAI222_X1 port map( A1 => n658, A2 => n803, B1 => n649, B2 => n676, 
                           C1 => n662, C2 => n673, ZN => n363);
   U340 : OAI222_X1 port map( A1 => n717, A2 => n319, B1 => n722, B2 => n366, 
                           C1 => n733, C2 => n332, ZN => n365);
   U341 : OAI222_X1 port map( A1 => n711, A2 => n319, B1 => n717, B2 => n366, 
                           C1 => n722, C2 => n332, ZN => n376);
   U342 : OAI222_X1 port map( A1 => n699, A2 => n319, B1 => n701, B2 => n366, 
                           C1 => n706, C2 => n332, ZN => n428);
   U343 : OAI222_X1 port map( A1 => n646, A2 => n685, B1 => n644, B2 => n799, 
                           C1 => n657, C2 => n673, ZN => n349);
   U344 : OAI222_X1 port map( A1 => n318, A2 => n319, B1 => n244, B2 => n757, 
                           C1 => n98, C2 => n672, ZN => n317);
   U345 : INV_X1 port map( A => n307, ZN => n757);
   U346 : OAI222_X1 port map( A1 => n658, A2 => n800, B1 => n649, B2 => n682, 
                           C1 => n662, C2 => n801, ZN => n312);
   U347 : OAI222_X1 port map( A1 => n659, A2 => n679, B1 => n649, B2 => n801, 
                           C1 => n663, C2 => n676, ZN => n339);
   U348 : OAI222_X1 port map( A1 => n659, A2 => n799, B1 => n649, B2 => n802, 
                           C1 => n663, C2 => n685, ZN => n262);
   U349 : NOR4_X1 port map( A1 => n444, A2 => n445, A3 => n446, A4 => n447, ZN 
                           => n443);
   U350 : OAI222_X1 port map( A1 => n659, A2 => n669, B1 => n649, B2 => n670, 
                           C1 => n663, C2 => n668, ZN => n447);
   U351 : OAI222_X1 port map( A1 => n722, A2 => n408, B1 => n733, B2 => n407, 
                           C1 => n716, C2 => n386, ZN => n438);
   U352 : OAI222_X1 port map( A1 => n660, A2 => n668, B1 => n649, B2 => n669, 
                           C1 => n661, C2 => n667, ZN => n466);
   U353 : NOR3_X1 port map( A1 => n410, A2 => n409, A3 => n411, ZN => n403);
   U354 : OAI22_X1 port map( A1 => n802, A2 => n249, B1 => n799, B2 => n247, ZN
                           => n411);
   U355 : OAI221_X1 port map( B1 => n695, B2 => n270, C1 => n691, C2 => n287, A
                           => n418, ZN => n409);
   U356 : OAI222_X1 port map( A1 => n717, A2 => n285, B1 => n347, B2 => n605, 
                           C1 => n712, C2 => n284, ZN => n345);
   U357 : NOR4_X1 port map( A1 => n348, A2 => n349, A3 => n350, A4 => n351, ZN 
                           => n347);
   U358 : OAI222_X1 port map( A1 => n660, A2 => n676, B1 => n649, B2 => n679, 
                           C1 => n661, C2 => n803, ZN => n351);
   U359 : OAI222_X1 port map( A1 => n697, A2 => n646, B1 => n699, B2 => n644, 
                           C1 => n655, C2 => n800, ZN => n274);
   U360 : OAI222_X1 port map( A1 => n646, A2 => n682, B1 => n644, B2 => n685, 
                           C1 => n656, C2 => n672, ZN => n361);
   U361 : OAI222_X1 port map( A1 => n646, A2 => n799, B1 => n644, B2 => n802, 
                           C1 => n655, C2 => n803, ZN => n337);
   U362 : OAI222_X1 port map( A1 => n646, A2 => n803, B1 => n644, B2 => n676, 
                           C1 => n656, C2 => n667, ZN => n445);
   U363 : OAI222_X1 port map( A1 => n646, A2 => n672, B1 => n644, B2 => n673, 
                           C1 => n656, C2 => n665, ZN => n493);
   U364 : OAI222_X1 port map( A1 => n646, A2 => n673, B1 => n644, B2 => n803, 
                           C1 => n655, C2 => n666, ZN => n464);
   U365 : OAI222_X1 port map( A1 => n699, A2 => n646, B1 => n701, B2 => n644, 
                           C1 => n656, C2 => n682, ZN => n260);
   U366 : OAI222_X1 port map( A1 => n646, A2 => n802, B1 => n691, B2 => n644, 
                           C1 => n657, C2 => n676, ZN => n323);
   U368 : OAI222_X1 port map( A1 => n702, A2 => n646, B1 => n707, B2 => n644, 
                           C1 => n657, C2 => n685, ZN => n251);
   U369 : OAI222_X1 port map( A1 => n703, A2 => n247, B1 => n321, B2 => n222, 
                           C1 => n706, C2 => n249, ZN => n320);
   U370 : NOR4_X1 port map( A1 => n322, A2 => n323, A3 => n324, A4 => n325, ZN 
                           => n321);
   U371 : OAI222_X1 port map( A1 => n659, A2 => n801, B1 => n649, B2 => n800, 
                           C1 => n663, C2 => n679, ZN => n325);
   U372 : OAI222_X1 port map( A1 => n722, A2 => n249, B1 => n716, B2 => n247, 
                           C1 => n272, C2 => n605, ZN => n267);
   U373 : NOR4_X1 port map( A1 => n273, A2 => n274, A3 => n275, A4 => n276, ZN 
                           => n272);
   U374 : OAI222_X1 port map( A1 => n660, A2 => n685, B1 => n649, B2 => n799, 
                           C1 => n661, C2 => n682, ZN => n276);
   U375 : AOI22_X1 port map( A1 => n609, A2 => n692, B1 => n624, B2 => n696, ZN
                           => n340);
   U376 : AOI22_X1 port map( A1 => n609, A2 => n710, B1 => n624, B2 => n715, ZN
                           => n263);
   U377 : AOI22_X1 port map( A1 => n609, A2 => n686, B1 => n624, B2 => n692, ZN
                           => n352);
   U378 : AOI22_X1 port map( A1 => n609, A2 => n704, B1 => n624, B2 => n710, ZN
                           => n277);
   U379 : AOI22_X1 port map( A1 => n609, A2 => n696, B1 => n624, B2 => n698, ZN
                           => n326);
   U380 : AOI22_X1 port map( A1 => n781, A2 => n698, B1 => n624, B2 => n700, ZN
                           => n313);
   U381 : AOI22_X1 port map( A1 => n609, A2 => n715, B1 => n624, B2 => n723, ZN
                           => n255);
   U382 : OAI222_X1 port map( A1 => n660, A2 => n682, B1 => n145, B2 => n685, 
                           C1 => n661, C2 => n800, ZN => n294);
   U383 : OAI222_X1 port map( A1 => n646, A2 => n679, B1 => n644, B2 => n801, 
                           C1 => n657, C2 => n669, ZN => n414);
   U384 : OAI222_X1 port map( A1 => n658, A2 => n671, B1 => n649, B2 => n672, 
                           C1 => n662, C2 => n670, ZN => n416);
   U385 : AOI221_X1 port map( B1 => n704, B2 => n789, C1 => n700, C2 => n794, A
                           => n178, ZN => n172);
   U386 : OAI22_X1 port map( A1 => n714, A2 => n649, B1 => n717, B2 => n642, ZN
                           => n178);
   U387 : OAI221_X1 port map( B1 => n784, B2 => n718, C1 => n722, C2 => n656, A
                           => n130, ZN => n124);
   U388 : AOI22_X1 port map( A1 => n789, A2 => n736, B1 => n794, B2 => n728, ZN
                           => n130);
   U389 : OAI221_X1 port map( B1 => n799, B2 => n270, C1 => n685, C2 => n287, A
                           => n468, ZN => n459);
   U390 : AOI222_X1 port map( A1 => n768, A2 => n698, B1 => n758, B2 => n696, 
                           C1 => n769, C2 => n693, ZN => n468);
   U391 : OAI221_X1 port map( B1 => n474, B2 => n334, C1 => n718, C2 => n407, A
                           => n475, ZN => n471);
   U393 : AOI22_X1 port map( A1 => n772, A2 => n723, B1 => n773, B2 => n710, ZN
                           => n475);
   U394 : NOR3_X1 port map( A1 => n485, A2 => n484, A3 => n486, ZN => n474);
   U395 : OAI22_X1 port map( A1 => n800, A2 => n249, B1 => n247, B2 => n801, ZN
                           => n486);
   U396 : OAI221_X1 port map( B1 => n697, B2 => n270, C1 => n695, C2 => n287, A
                           => n392, ZN => n390);
   U397 : AOI222_X1 port map( A1 => n768, A2 => r1(28), B1 => n758, B2 => n710,
                           C1 => n769, C2 => n704, ZN => n392);
   U398 : OAI221_X1 port map( B1 => n457, B2 => n334, C1 => n722, C2 => n407, A
                           => n458, ZN => n452);
   U399 : AOI22_X1 port map( A1 => n772, A2 => n727, B1 => n773, B2 => n715, ZN
                           => n458);
   U400 : NOR3_X1 port map( A1 => n459, A2 => n460, A3 => n461, ZN => n457);
   U401 : OAI22_X1 port map( A1 => n682, A2 => n249, B1 => n247, B2 => n800, ZN
                           => n461);
   U402 : OAI221_X1 port map( B1 => n706, B2 => n270, C1 => n702, C2 => n287, A
                           => n353, ZN => n344);
   U403 : AOI222_X1 port map( A1 => n768, A2 => n736, B1 => n758, B2 => n729, 
                           C1 => n769, C2 => n724, ZN => n353);
   U404 : AOI22_X1 port map( A1 => n781, A2 => n700, B1 => n624, B2 => n704, ZN
                           => n295);
   U405 : OAI221_X1 port map( B1 => n784, B2 => n699, C1 => n655, C2 => n702, A
                           => n167, ZN => n164);
   U406 : AOI22_X1 port map( A1 => n793, A2 => n727, B1 => n787, B2 => n736, ZN
                           => n167);
   U407 : NOR3_X1 port map( A1 => n119, A2 => n582, A3 => n158, ZN => n125);
   U409 : OAI21_X1 port map( B1 => n371, B2 => n297, A => n386, ZN => n385);
   U410 : OAI211_X1 port map( C1 => n722, C2 => n287, A => n271, B => n289, ZN 
                           => n279);
   U411 : OAI221_X1 port map( B1 => n98, B2 => n666, C1 => n101, C2 => n667, A 
                           => n400, ZN => N2064);
   U412 : OAI21_X1 port map( B1 => n401, B2 => n402, A => n123, ZN => n400);
   U413 : OAI222_X1 port map( A1 => n722, A2 => n372, B1 => n733, B2 => n386, 
                           C1 => n716, C2 => n387, ZN => n402);
   U414 : OAI221_X1 port map( B1 => n750, B2 => n403, C1 => n297, C2 => n404, A
                           => n405, ZN => n401);
   U415 : AOI221_X1 port map( B1 => n134, B2 => n299, C1 => n300, C2 => n282, A
                           => n162, ZN => n298);
   U416 : AOI21_X1 port map( B1 => n301, B2 => n302, A => n753, ZN => n300);
   U417 : OAI221_X1 port map( B1 => n98, B2 => n799, C1 => n101, C2 => n802, A 
                           => n191, ZN => N2079);
   U418 : AOI221_X1 port map( B1 => n128, B2 => n192, C1 => n193, C2 => n777, A
                           => n162, ZN => n191);
   U419 : INV_X1 port map( A => n194, ZN => n777);
   U420 : OAI21_X1 port map( B1 => n200, B2 => n566, A => n163, ZN => n192);
   U421 : OAI221_X1 port map( B1 => n98, B2 => n722, C1 => n733, C2 => n101, A 
                           => n103, ZN => N2089);
   U422 : OAI21_X1 port map( B1 => n104, B2 => n752, A => n776, ZN => n103);
   U423 : OAI221_X1 port map( B1 => n733, B2 => n660, C1 => n722, C2 => n661, A
                           => n139, ZN => n135);
   U424 : OAI22_X1 port map( A1 => n788, A2 => n711, B1 => n655, B2 => n716, ZN
                           => n140);
   U425 : NOR2_X1 port map( A1 => n158, A2 => n775, ZN => n186);
   U426 : OAI22_X1 port map( A1 => n658, A2 => n699, B1 => n649, B2 => n701, ZN
                           => n206);
   U427 : OAI22_X1 port map( A1 => n708, A2 => n145, B1 => n714, B2 => n642, ZN
                           => n190);
   U428 : OAI22_X1 port map( A1 => n98, A2 => n665, B1 => n318, B2 => n407, ZN 
                           => n422);
   U429 : OAI221_X1 port map( B1 => n743, B2 => n159, C1 => n98, C2 => n695, A 
                           => n160, ZN => N2082);
   U430 : NOR2_X1 port map( A1 => n164, A2 => n165, ZN => n159);
   U431 : AOI21_X1 port map( B1 => n696, B2 => n601, A => n749, ZN => n160);
   U432 : OAI221_X1 port map( B1 => n722, B2 => n642, C1 => n719, C2 => n145, A
                           => n166, ZN => n165);
   U433 : OAI221_X1 port map( B1 => n747, B2 => n341, C1 => n98, C2 => n670, A 
                           => n342, ZN => N2068);
   U434 : AOI21_X1 port map( B1 => r1(9), B2 => n601, A => n748, ZN => n342);
   U435 : NOR3_X1 port map( A1 => n344, A2 => n345, A3 => n346, ZN => n341);
   U436 : OAI22_X1 port map( A1 => n699, A2 => n249, B1 => n697, B2 => n247, ZN
                           => n346);
   U437 : AOI22_X1 port map( A1 => n779, A2 => n716, B1 => n232, B2 => n644, ZN
                           => n231);
   U438 : OAI22_X1 port map( A1 => r1(27), A2 => n646, B1 => n233, B2 => n234, 
                           ZN => n232);
   U439 : OAI221_X1 port map( B1 => n659, B2 => n695, C1 => n663, C2 => n691, A
                           => n236, ZN => n233);
   U440 : OAI21_X1 port map( B1 => n334, B2 => n297, A => n158, ZN => n391);
   U441 : INV_X1 port map( A => n713, ZN => n710);
   U442 : INV_X1 port map( A => n707, ZN => n704);
   U443 : OAI22_X1 port map( A1 => n722, A2 => n145, B1 => n574, B2 => n154, ZN
                           => n152);
   U444 : AOI22_X1 port map( A1 => n155, A2 => n658, B1 => n789, B2 => n715, ZN
                           => n154);
   U445 : OAI221_X1 port map( B1 => n655, B2 => n708, C1 => n662, C2 => n713, A
                           => n156, ZN => n155);
   U446 : OAI22_X1 port map( A1 => n782, A2 => n779, B1 => n644, B2 => n724, ZN
                           => n216);
   U447 : INV_X1 port map( A => n217, ZN => n782);
   U448 : OAI22_X1 port map( A1 => r1(28), A2 => n646, B1 => n218, B2 => n219, 
                           ZN => n217);
   U449 : INV_X1 port map( A => n681, ZN => n682);
   U450 : INV_X1 port map( A => r2(3), ZN => n795);
   U451 : OAI211_X1 port map( C1 => n101, C2 => n685, A => n223, B => n224, ZN 
                           => N2077);
   U452 : AOI221_X1 port map( B1 => n226, B2 => n227, C1 => n609, C2 => n733, A
                           => n228, ZN => n225);
   U453 : OAI211_X1 port map( C1 => n101, C2 => n801, A => n742, B => n256, ZN 
                           => N2074);
   U454 : OAI222_X1 port map( A1 => n722, A2 => n247, B1 => n258, B2 => n222, 
                           C1 => n733, C2 => n249, ZN => n257);
   U455 : NOR4_X1 port map( A1 => n259, A2 => n260, A3 => n261, A4 => n262, ZN 
                           => n258);
   U456 : OAI211_X1 port map( C1 => n101, C2 => n699, A => n141, B => n148, ZN 
                           => N2083);
   U457 : NOR3_X1 port map( A1 => n150, A2 => n144, A3 => n151, ZN => n149);
   U458 : OAI211_X1 port map( C1 => n101, C2 => n799, A => n208, B => n209, ZN 
                           => N2078);
   U459 : AOI221_X1 port map( B1 => n210, B2 => n193, C1 => n609, C2 => n776, A
                           => n162, ZN => n209);
   U460 : OAI211_X1 port map( C1 => n202, C2 => n740, A => n213, B => n163, ZN 
                           => n212);
   U461 : NOR4_X1 port map( A1 => n505, A2 => r2(30), A3 => r2(5), A4 => r2(31)
                           , ZN => n504);
   U462 : NOR4_X1 port map( A1 => n508, A2 => r2(10), A3 => r2(12), A4 => 
                           r2(11), ZN => n501);
   U463 : NAND2_X1 port map( A1 => n737, A2 => n752, ZN => n100);
   U464 : AOI22_X1 port map( A1 => n790, A2 => n686, B1 => n760, B2 => n692, ZN
                           => n373);
   U465 : AOI221_X1 port map( B1 => n755, B2 => n698, C1 => n767, C2 => n696, A
                           => n376, ZN => n375);
   U466 : BUF_X1 port map( A => r1(22), Z => n692);
   U467 : BUF_X1 port map( A => r1(22), Z => n693);
   U468 : BUF_X1 port map( A => n720, Z => n723);
   U469 : BUF_X1 port map( A => n720, Z => n724);
   U470 : BUF_X1 port map( A => n721, Z => n726);
   U471 : BUF_X1 port map( A => r1(18), Z => n683);
   U472 : OR3_X1 port map( A1 => r2(15), A2 => r2(14), A3 => r2(13), ZN => n508
                           );
   U473 : BUF_X1 port map( A => n721, Z => n725);
   U474 : BUF_X1 port map( A => r1(18), Z => n684);
   U475 : AOI222_X1 port map( A1 => n771, A2 => n715, B1 => n773, B2 => n729, 
                           C1 => n765, C2 => n725, ZN => n420);
   U476 : AOI211_X1 port map( C1 => r1(4), C2 => n601, A => n422, B => n423, ZN
                           => n421);
   U477 : AOI22_X1 port map( A1 => n762, A2 => n710, B1 => n424, B2 => n268, ZN
                           => n419);
   U478 : BUF_X1 port map( A => r1(14), Z => n677);
   U479 : OR3_X1 port map( A1 => n158, A2 => n775, A3 => n605, ZN => n211);
   U480 : BUF_X1 port map( A => r1(13), Z => n674);
   U481 : BUF_X1 port map( A => r1(22), Z => n694);
   U482 : BUF_X1 port map( A => r1(14), Z => n678);
   U483 : BUF_X1 port map( A => r1(13), Z => n675);
   U484 : BUF_X1 port map( A => r1(30), Z => n731);
   U485 : BUF_X1 port map( A => r1(30), Z => n732);
   U486 : AOI22_X1 port map( A1 => n680, A2 => n781, B1 => n624, B2 => n683, ZN
                           => n417);
   U487 : AOI22_X1 port map( A1 => n674, A2 => n781, B1 => n678, B2 => n624, ZN
                           => n496);
   U488 : INV_X1 port map( A => r1(19), ZN => n799);
   U489 : INV_X1 port map( A => r1(20), ZN => n802);
   U490 : INV_X1 port map( A => r1(16), ZN => n800);
   U491 : AOI221_X1 port map( B1 => n778, B2 => n684, C1 => r1(19), C2 => n788,
                           A => n243, ZN => n242);
   U492 : OAI22_X1 port map( A1 => n662, A2 => n802, B1 => n658, B2 => n691, ZN
                           => n243);
   U493 : AOI221_X1 port map( B1 => r1(5), B2 => n778, C1 => r1(15), C2 => n792
                           , A => n434, ZN => n433);
   U494 : OAI22_X1 port map( A1 => n230, A2 => n682, B1 => n227, B2 => n800, ZN
                           => n434);
   U495 : OAI22_X1 port map( A1 => n799, A2 => n230, B1 => n227, B2 => n685, ZN
                           => n399);
   U496 : INV_X1 port map( A => r1(15), ZN => n801);
   U497 : INV_X1 port map( A => r1(12), ZN => n803);
   U498 : OAI221_X1 port map( B1 => n659, B2 => n697, C1 => n663, C2 => n695, A
                           => n221, ZN => n218);
   U499 : OAI221_X1 port map( B1 => n454, B2 => n469, C1 => n318, C2 => n105, A
                           => n470, ZN => N2060);
   U500 : NOR2_X1 port map( A1 => n471, A2 => n472, ZN => n469);
   U501 : OAI221_X1 port map( B1 => n705, B2 => n386, C1 => n733, C2 => n455, A
                           => n473, ZN => n472);
   U502 : AOI21_X1 port map( B1 => n356, B2 => n357, A => n747, ZN => n355);
   U503 : AOI221_X1 port map( B1 => n755, B2 => n700, C1 => n767, C2 => n698, A
                           => n365, ZN => n356);
   U504 : OAI211_X1 port map( C1 => n101, C2 => n669, A => n367, B => n368, ZN 
                           => N2066);
   U505 : OAI21_X1 port map( B1 => n371, B2 => n620, A => n372, ZN => n370);
   U506 : OAI211_X1 port map( C1 => n101, C2 => n800, A => n742, B => n245, ZN 
                           => N2075);
   U507 : OAI222_X1 port map( A1 => n733, A2 => n247, B1 => n248, B2 => n222, 
                           C1 => n738, C2 => n249, ZN => n246);
   U508 : NOR4_X1 port map( A1 => n250, A2 => n251, A3 => n252, A4 => n253, ZN 
                           => n248);
   U509 : OAI211_X1 port map( C1 => n101, C2 => n682, A => n223, B => n237, ZN 
                           => N2076);
   U510 : NAND4_X1 port map( A1 => n239, A2 => n240, A3 => n241, A4 => n242, ZN
                           => n238);
   U511 : NAND4_X1 port map( A1 => n378, A2 => n379, A3 => n380, A4 => n381, ZN
                           => n377);
   U512 : AOI222_X1 port map( A1 => r1(10), A2 => n794, B1 => r1(12), B2 => 
                           n574, C1 => r1(11), C2 => n789, ZN => n378);
   U513 : AOI222_X1 port map( A1 => r1(9), A2 => n788, B1 => n681, B2 => n779, 
                           C1 => r1(16), C2 => n791, ZN => n380);
   U514 : NAND4_X1 port map( A1 => n430, A2 => n431, A3 => n432, A4 => n433, ZN
                           => n429);
   U515 : AOI222_X1 port map( A1 => r1(7), A2 => n794, B1 => r1(9), B2 => n574,
                           C1 => r1(8), C2 => n789, ZN => n430);
   U516 : AOI222_X1 port map( A1 => r1(6), A2 => n788, B1 => n677, B2 => n779, 
                           C1 => n675, C2 => n791, ZN => n432);
   U517 : AOI222_X1 port map( A1 => r1(9), A2 => n794, B1 => r1(11), B2 => n625
                           , C1 => r1(10), C2 => n789, ZN => n395);
   U518 : AOI222_X1 port map( A1 => r1(8), A2 => n788, B1 => r1(16), B2 => n779
                           , C1 => r1(15), C2 => n791, ZN => n397);
   U519 : NAND4_X1 port map( A1 => n327, A2 => n328, A3 => n329, A4 => n330, ZN
                           => N2069);
   U520 : AOI222_X1 port map( A1 => n769, A2 => n730, B1 => n759, B2 => n723, 
                           C1 => n770, C2 => n715, ZN => n330);
   U521 : AOI21_X1 port map( B1 => r1(10), B2 => n601, A => n748, ZN => n327);
   U522 : AOI221_X1 port map( B1 => n755, B2 => n710, C1 => n767, C2 => n704, A
                           => n331, ZN => n329);
   U523 : AOI21_X1 port map( B1 => n440, B2 => n441, A => n747, ZN => n439);
   U532 : AOI221_X1 port map( B1 => n755, B2 => r1(20), C1 => n767, C2 => 
                           r1(19), A => n449, ZN => n440);
   U541 : OAI222_X1 port map( A1 => n697, A2 => n319, B1 => n699, B2 => n366, 
                           C1 => n702, C2 => n332, ZN => n449);
   U542 : AOI22_X1 port map( A1 => n790, A2 => n683, B1 => n760, B2 => r1(19), 
                           ZN => n425);
   U543 : AOI221_X1 port map( B1 => n755, B2 => n690, C1 => n767, C2 => r1(20),
                           A => n428, ZN => n427);
   U544 : AOI222_X1 port map( A1 => n770, A2 => n693, B1 => n214, B2 => n429, 
                           C1 => n759, C2 => n696, ZN => n426);
   U545 : INV_X1 port map( A => r1(23), ZN => n697);
   U546 : AOI222_X1 port map( A1 => n755, A2 => n715, B1 => n759, B2 => n729, 
                           C1 => n770, C2 => n725, ZN => n315);
   U547 : AOI211_X1 port map( C1 => r1(11), C2 => n601, A => n317, B => n748, 
                           ZN => n316);
   U548 : AOI22_X1 port map( A1 => n767, A2 => n710, B1 => n320, B2 => n745, ZN
                           => n314);
   U549 : BUF_X1 port map( A => r1(17), Z => n680);
   U550 : AOI22_X1 port map( A1 => n779, A2 => n736, B1 => n791, B2 => n728, ZN
                           => n179);
   U551 : AOI22_X1 port map( A1 => n182, A2 => n118, B1 => n183, B2 => n157, ZN
                           => n180);
   U552 : AOI221_X1 port map( B1 => n771, B2 => r1(27), C1 => n762, C2 => n704,
                           A => n438, ZN => n437);
   U553 : AOI21_X1 port map( B1 => r1(3), B2 => n601, A => n423, ZN => n435);
   U554 : BUF_X1 port map( A => r1(17), Z => n681);
   U555 : OAI21_X1 port map( B1 => n452, B2 => n453, A => n766, ZN => n450);
   U556 : OAI221_X1 port map( B1 => n711, B2 => n386, C1 => n740, C2 => n455, A
                           => n456, ZN => n453);
   U557 : BUF_X1 port map( A => r1(29), Z => n720);
   U558 : BUF_X1 port map( A => r1(29), Z => n721);
   U559 : AOI22_X1 port map( A1 => n609, A2 => r1(20), B1 => n624, B2 => n687, 
                           ZN => n364);
   U560 : AOI22_X1 port map( A1 => r1(15), A2 => n781, B1 => r1(16), B2 => n624
                           , ZN => n448);
   U561 : AOI22_X1 port map( A1 => n677, A2 => n609, B1 => r1(15), B2 => n624, 
                           ZN => n467);
   U562 : INV_X1 port map( A => log, ZN => n752);
   U563 : NAND2_X1 port map( A1 => n499, A2 => n490, ZN => n153);
   U564 : OAI211_X1 port map( C1 => n101, C2 => n670, A => n343, B => n354, ZN 
                           => N2067);
   U565 : AOI22_X1 port map( A1 => n152, A2 => n642, B1 => n786, B2 => n728, ZN
                           => n151);
   U566 : AOI222_X1 port map( A1 => n693, A2 => n574, B1 => n793, B2 => n698, 
                           C1 => n696, C2 => n786, ZN => n241);
   U567 : AOI222_X1 port map( A1 => r1(10), A2 => n786, B1 => r1(11), B2 => 
                           n793, C1 => r1(12), C2 => n787, ZN => n431);
   U568 : AOI222_X1 port map( A1 => n674, A2 => n786, B1 => n677, B2 => n793, 
                           C1 => r1(15), C2 => n787, ZN => n379);
   U569 : AOI222_X1 port map( A1 => r1(12), A2 => n786, B1 => n674, B2 => n793,
                           C1 => n678, C2 => n787, ZN => n396);
   U570 : AOI22_X1 port map( A1 => n698, A2 => n786, B1 => n696, B2 => n574, ZN
                           => n235);
   U571 : AOI22_X1 port map( A1 => n786, A2 => n700, B1 => n698, B2 => n574, ZN
                           => n220);
   U572 : CLKBUF_X1 port map( A => n197, Z => n643);
   U573 : NAND2_X1 port map( A1 => n478, A2 => n651, ZN => n197);
   U574 : OAI22_X1 port map( A1 => n195, A2 => n792, B1 => n196, B2 => n736, ZN
                           => n194);
   U575 : OAI22_X1 port map( A1 => n726, A2 => n196, B1 => n792, B2 => n231, ZN
                           => n226);
   U576 : AOI22_X1 port map( A1 => n733, A2 => n792, B1 => n196, B2 => n216, ZN
                           => n210);
   U577 : OAI221_X1 port map( B1 => n654, B2 => n803, C1 => n695, C2 => n196, A
                           => n326, ZN => n322);
   U578 : OAI221_X1 port map( B1 => n682, B2 => n654, C1 => n711, C2 => n196, A
                           => n255, ZN => n250);
   U579 : OAI221_X1 port map( B1 => n654, B2 => n801, C1 => n702, C2 => n196, A
                           => n277, ZN => n273);
   U580 : OAI221_X1 port map( B1 => n654, B2 => n672, C1 => n802, C2 => n196, A
                           => n352, ZN => n348);
   U581 : AOI21_X1 port map( B1 => n196, B2 => n202, A => n739, ZN => n183);
   U582 : OAI221_X1 port map( B1 => n654, B2 => n800, C1 => n709, C2 => n196, A
                           => n263, ZN => n259);
   U583 : OAI221_X1 port map( B1 => n654, B2 => n673, C1 => n691, C2 => n196, A
                           => n340, ZN => n336);
   U584 : OAI221_X1 port map( B1 => n654, B2 => n676, C1 => n697, C2 => n196, A
                           => n313, ZN => n309);
   U585 : OAI221_X1 port map( B1 => n573, B2 => n679, C1 => n699, C2 => n196, A
                           => n295, ZN => n291);
   U587 : AOI22_X1 port map( A1 => r1(1), A2 => n600, B1 => r1(2), B2 => n601, 
                           ZN => n451);
   U588 : OR3_X1 port map( A1 => n648, A2 => n600, A3 => n100, ZN => n102);
   U589 : AOI22_X1 port map( A1 => r1(0), A2 => n600, B1 => r1(1), B2 => n601, 
                           ZN => n470);
   U590 : AOI22_X1 port map( A1 => r1(26), A2 => n600, B1 => r1(27), B2 => n601
                           , ZN => n122);
   U591 : AOI22_X1 port map( A1 => n246, A2 => n745, B1 => r1(15), B2 => n600, 
                           ZN => n245);
   U592 : AOI22_X1 port map( A1 => n143, A2 => n746, B1 => n698, B2 => n600, ZN
                           => n142);
   U593 : AOI22_X1 port map( A1 => n767, A2 => n727, B1 => n674, B2 => n600, ZN
                           => n265);
   U594 : AOI22_X1 port map( A1 => n762, A2 => n727, B1 => r1(6), B2 => n600, 
                           ZN => n367);
   U595 : AOI22_X1 port map( A1 => n134, A2 => n212, B1 => n684, B2 => n600, ZN
                           => n208);
   U596 : AOI221_X1 port map( B1 => r1(20), B2 => n600, C1 => n689, C2 => n601,
                           A => n116, ZN => n181);
   U597 : AOI221_X1 port map( B1 => r1(2), B2 => n600, C1 => n772, C2 => n776, 
                           A => n439, ZN => n436);
   U598 : AOI222_X1 port map( A1 => n677, A2 => n600, B1 => n745, B2 => n257, 
                           C1 => n767, C2 => n736, ZN => n256);
   U599 : AOI222_X1 port map( A1 => r1(16), A2 => n600, B1 => n229, B2 => n238,
                           C1 => n790, C2 => n776, ZN => n237);
   U600 : AOI221_X1 port map( B1 => n688, B2 => n600, C1 => n694, C2 => n601, A
                           => n116, ZN => n170);
   U601 : AOI221_X1 port map( B1 => n710, B2 => n600, C1 => r1(28), C2 => n601,
                           A => n116, ZN => n115);
   U602 : AOI221_X1 port map( B1 => n696, B2 => n600, C1 => n793, C2 => n776, A
                           => n149, ZN => n148);
   U603 : AOI222_X1 port map( A1 => n704, A2 => n601, B1 => n134, B2 => n579, 
                           C1 => r1(25), C2 => n600, ZN => n133);
   U604 : NOR4_X1 port map( A1 => n297, A2 => n648, A3 => n601, A4 => n600, ZN 
                           => n128);
   U605 : BUF_X1 port map( A => n99, Z => n647);
   U606 : AOI22_X1 port map( A1 => n111, A2 => n107, B1 => n112, B2 => n784, ZN
                           => n109);
   U607 : AND4_X1 port map( A1 => n105, A2 => n761, A3 => n106, A4 => n107, ZN 
                           => n104);
   U608 : AOI22_X1 port map( A1 => n693, A2 => n107, B1 => n696, B2 => n788, ZN
                           => n188);
   U609 : AOI22_X1 port map( A1 => r1(26), A2 => n107, B1 => n786, B2 => n736, 
                           ZN => n146);
   U610 : AOI221_X1 port map( B1 => n696, B2 => n107, C1 => n698, C2 => n788, A
                           => n175, ZN => n173);
   U611 : INV_X1 port map( A => n107, ZN => n784);
   U612 : AOI22_X1 port map( A1 => n689, A2 => n107, B1 => n786, B2 => n704, ZN
                           => n203);
   U613 : CLKBUF_X1 port map( A => n168, Z => n645);
   U614 : NAND2_X1 port map( A1 => n478, A2 => n653, ZN => n168);
   U615 : NAND2_X1 port map( A1 => n478, A2 => n481, ZN => n408);
   U616 : NAND2_X1 port map( A1 => n481, A2 => n491, ZN => n287);
   U617 : NAND2_X1 port map( A1 => n481, A2 => n499, ZN => n332);
   U618 : NAND2_X1 port map( A1 => n481, A2 => n497, ZN => n319);
   U619 : NAND2_X1 port map( A1 => n482, A2 => n481, ZN => n476);
   U620 : OAI22_X1 port map( A1 => n733, A2 => n607, B1 => n722, B2 => n640, ZN
                           => n175);
   U621 : OAI222_X1 port map( A1 => n607, A2 => n799, B1 => n640, B2 => n685, 
                           C1 => n642, C2 => n682, ZN => n324);
   U622 : OAI222_X1 port map( A1 => n699, A2 => n607, B1 => n640, B2 => n697, 
                           C1 => n642, C2 => n695, ZN => n252);
   U623 : OAI222_X1 port map( A1 => n607, A2 => n695, B1 => n640, B2 => n691, 
                           C1 => n642, C2 => n802, ZN => n275);
   U624 : OAI222_X1 port map( A1 => n607, A2 => n682, B1 => n640, B2 => n800, 
                           C1 => n642, C2 => n801, ZN => n350);
   U625 : OAI222_X1 port map( A1 => n697, A2 => n607, B1 => n640, B2 => n695, 
                           C1 => n642, C2 => n691, ZN => n261);
   U626 : OAI222_X1 port map( A1 => n607, A2 => n685, B1 => n640, B2 => n682, 
                           C1 => n642, C2 => n800, ZN => n338);
   U627 : OAI222_X1 port map( A1 => n607, A2 => n672, B1 => n640, B2 => n671, 
                           C1 => n642, C2 => n670, ZN => n465);
   U628 : OAI221_X1 port map( B1 => n702, B2 => n640, C1 => n709, C2 => n607, A
                           => n235, ZN => n234);
   U629 : OAI222_X1 port map( A1 => n607, A2 => n671, B1 => n640, B2 => n670, 
                           C1 => n642, C2 => n669, ZN => n494);
   U630 : OAI222_X1 port map( A1 => n607, A2 => n676, B1 => n640, B2 => n803, 
                           C1 => n642, C2 => n673, ZN => n415);
   U631 : OAI221_X1 port map( B1 => n705, B2 => n640, C1 => n714, C2 => n607, A
                           => n220, ZN => n219);
   U632 : OAI222_X1 port map( A1 => n607, A2 => n673, B1 => n640, B2 => n672, 
                           C1 => n642, C2 => n671, ZN => n446);
   U633 : OAI222_X1 port map( A1 => n607, A2 => n802, B1 => n640, B2 => n799, 
                           C1 => n642, C2 => n685, ZN => n311);
   U634 : OAI222_X1 port map( A1 => n607, A2 => n800, B1 => n640, B2 => n801, 
                           C1 => n642, C2 => n679, ZN => n362);
   U635 : OAI222_X1 port map( A1 => n607, A2 => n691, B1 => n640, B2 => n802, 
                           C1 => n642, C2 => n799, ZN => n293);
   U636 : INV_X1 port map( A => n177, ZN => n793);
   U637 : NAND2_X1 port map( A1 => n176, A2 => n177, ZN => n150);
   U638 : NAND4_X1 port map( A1 => n504, A2 => n501, A3 => n503, A4 => n502, ZN
                           => n99);
   U639 : AND4_X2 port map( A1 => n136, A2 => n108, A3 => n137, A4 => n138, ZN 
                           => n107);
   U640 : INV_X1 port map( A => n626, ZN => n785);
   U641 : NAND2_X1 port map( A1 => n489, A2 => n606, ZN => n108);
   U642 : NAND2_X1 port map( A1 => n497, A2 => n651, ZN => n137);
   U643 : NAND2_X1 port map( A1 => n497, A2 => n652, ZN => n138);
   U644 : AOI22_X1 port map( A1 => n574, A2 => n776, B1 => n112, B2 => n785, ZN
                           => n132);
   U645 : NAND2_X1 port map( A1 => n737, A2 => n785, ZN => n129);
   U646 : NOR3_X1 port map( A1 => n119, A2 => n789, A3 => n785, ZN => n113);
   U647 : AOI221_X1 port map( B1 => r1(8), B2 => n778, C1 => n683, C2 => n792, 
                           A => n382, ZN => n381);
   U648 : INV_X1 port map( A => n573, ZN => n778);
   U649 : NOR3_X1 port map( A1 => n786, A2 => n625, A3 => n150, ZN => n136);
   U650 : AOI211_X1 port map( C1 => n128, C2 => n279, A => n162, B => n280, ZN 
                           => n278);
   U651 : INV_X1 port map( A => r2(0), ZN => n798);
   U652 : OAI21_X1 port map( B1 => n389, B2 => n390, A => n391, ZN => n388);
   U653 : INV_X1 port map( A => r1(2), ZN => n664);
   U654 : INV_X1 port map( A => r1(3), ZN => n665);
   U655 : INV_X1 port map( A => r1(4), ZN => n666);
   U656 : INV_X1 port map( A => r1(5), ZN => n667);
   U657 : INV_X1 port map( A => r1(6), ZN => n668);
   U658 : INV_X1 port map( A => r1(7), ZN => n669);
   U659 : INV_X1 port map( A => r1(8), ZN => n670);
   U660 : INV_X1 port map( A => r1(9), ZN => n671);
   U661 : INV_X1 port map( A => r1(10), ZN => n672);
   U662 : INV_X1 port map( A => r1(11), ZN => n673);
   U663 : CLKBUF_X1 port map( A => r1(21), Z => n686);
   U664 : CLKBUF_X1 port map( A => r1(21), Z => n687);
   U665 : CLKBUF_X1 port map( A => r1(21), Z => n688);
   U666 : CLKBUF_X1 port map( A => r1(21), Z => n689);
   U667 : CLKBUF_X1 port map( A => r1(21), Z => n690);
   U668 : INV_X1 port map( A => n697, ZN => n696);
   U669 : INV_X1 port map( A => n699, ZN => n698);
   U670 : INV_X1 port map( A => r1(25), ZN => n701);
   U671 : INV_X1 port map( A => r1(25), ZN => n702);
   U672 : INV_X1 port map( A => r1(25), ZN => n703);
   U673 : INV_X1 port map( A => r1(26), ZN => n705);
   U674 : INV_X1 port map( A => r1(26), ZN => n706);
   U675 : INV_X1 port map( A => r1(26), ZN => n707);
   U676 : INV_X1 port map( A => r1(26), ZN => n708);
   U677 : INV_X1 port map( A => r1(26), ZN => n709);
   U678 : INV_X1 port map( A => r1(27), ZN => n711);
   U679 : INV_X1 port map( A => r1(27), ZN => n712);
   U680 : INV_X1 port map( A => r1(27), ZN => n713);
   U681 : INV_X1 port map( A => r1(27), ZN => n714);
   U682 : INV_X1 port map( A => r1(28), ZN => n716);
   U683 : INV_X1 port map( A => r1(28), ZN => n717);
   U684 : INV_X1 port map( A => r1(28), ZN => n718);
   U685 : INV_X1 port map( A => r1(28), ZN => n719);
   U686 : CLKBUF_X1 port map( A => r1(31), Z => n734);
   U687 : CLKBUF_X1 port map( A => r1(31), Z => n735);
   U688 : INV_X1 port map( A => n741, ZN => n737);
   U689 : INV_X1 port map( A => n734, ZN => n738);
   U690 : INV_X1 port map( A => n735, ZN => n739);
   U691 : INV_X1 port map( A => n735, ZN => n740);
   U692 : INV_X1 port map( A => r1(31), ZN => n741);
   U693 : INV_X2 port map( A => n270, ZN => n755);
   U694 : INV_X2 port map( A => n287, ZN => n767);
   U695 : INV_X2 port map( A => n153, ZN => n786);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity shifter_sx_nbit32 is

   port( r1, r2 : in std_logic_vector (31 downto 0);  data_out : out 
         std_logic_vector (31 downto 0));

end shifter_sx_nbit32;

architecture SYN_beh of shifter_sx_nbit32 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N1155, N1156, N1157, N1158, N1159, N1160, N1162, N1163, N1164, N1165,
      N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, 
      N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, n1,
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n451, n452, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677 : 
      std_logic;

begin
   
   data_out_reg_31_inst : DLH_X1 port map( G => n1, D => n629, Q => 
                           data_out(31));
   data_out_reg_30_inst : DLH_X1 port map( G => n1, D => N1185, Q => 
                           data_out(30));
   data_out_reg_29_inst : DLH_X1 port map( G => n1, D => N1184, Q => 
                           data_out(29));
   data_out_reg_28_inst : DLH_X1 port map( G => n1, D => N1183, Q => 
                           data_out(28));
   data_out_reg_27_inst : DLH_X1 port map( G => n1, D => N1182, Q => 
                           data_out(27));
   data_out_reg_26_inst : DLH_X1 port map( G => n1, D => N1181, Q => 
                           data_out(26));
   data_out_reg_25_inst : DLH_X1 port map( G => n1, D => N1180, Q => 
                           data_out(25));
   data_out_reg_24_inst : DLH_X1 port map( G => n1, D => N1179, Q => 
                           data_out(24));
   data_out_reg_23_inst : DLH_X1 port map( G => n1, D => N1178, Q => 
                           data_out(23));
   data_out_reg_22_inst : DLH_X1 port map( G => n1, D => N1177, Q => 
                           data_out(22));
   data_out_reg_21_inst : DLH_X1 port map( G => n1, D => N1176, Q => 
                           data_out(21));
   data_out_reg_20_inst : DLH_X1 port map( G => n1, D => N1175, Q => 
                           data_out(20));
   data_out_reg_19_inst : DLH_X1 port map( G => n1, D => N1174, Q => 
                           data_out(19));
   data_out_reg_18_inst : DLH_X1 port map( G => n1, D => N1173, Q => 
                           data_out(18));
   data_out_reg_17_inst : DLH_X1 port map( G => n1, D => N1172, Q => 
                           data_out(17));
   data_out_reg_16_inst : DLH_X1 port map( G => n1, D => N1171, Q => 
                           data_out(16));
   data_out_reg_15_inst : DLH_X1 port map( G => n1, D => N1170, Q => 
                           data_out(15));
   data_out_reg_14_inst : DLH_X1 port map( G => n1, D => N1169, Q => 
                           data_out(14));
   data_out_reg_13_inst : DLH_X1 port map( G => n1, D => N1168, Q => 
                           data_out(13));
   data_out_reg_12_inst : DLH_X1 port map( G => n1, D => N1167, Q => 
                           data_out(12));
   data_out_reg_11_inst : DLH_X1 port map( G => n1, D => N1166, Q => 
                           data_out(11));
   data_out_reg_10_inst : DLH_X1 port map( G => n1, D => N1165, Q => 
                           data_out(10));
   data_out_reg_9_inst : DLH_X1 port map( G => n1, D => N1164, Q => data_out(9)
                           );
   data_out_reg_8_inst : DLH_X1 port map( G => n1, D => N1163, Q => data_out(8)
                           );
   data_out_reg_7_inst : DLH_X1 port map( G => n1, D => N1162, Q => data_out(7)
                           );
   data_out_reg_6_inst : DLH_X1 port map( G => n1, D => n452, Q => data_out(6))
                           ;
   data_out_reg_5_inst : DLH_X1 port map( G => n1, D => N1160, Q => data_out(5)
                           );
   data_out_reg_4_inst : DLH_X1 port map( G => n1, D => N1159, Q => data_out(4)
                           );
   data_out_reg_3_inst : DLH_X1 port map( G => n1, D => N1158, Q => data_out(3)
                           );
   data_out_reg_2_inst : DLH_X1 port map( G => n1, D => N1157, Q => data_out(2)
                           );
   data_out_reg_1_inst : DLH_X1 port map( G => n1, D => N1156, Q => data_out(1)
                           );
   data_out_reg_0_inst : DLH_X1 port map( G => n1, D => N1155, Q => data_out(0)
                           );
   n1 <= '1';
   U349 : OR4_X2 port map( A1 => n87, A2 => n93, A3 => n664, A4 => n657, ZN => 
                           n153);
   U367 : NAND2_X2 port map( A1 => n440, A2 => n433, ZN => n167);
   U476 : OAI33_X1 port map( A1 => n557, A2 => n85, A3 => n86, B1 => n88, B2 =>
                           n87, B3 => n89, ZN => n84);
   U477 : NAND3_X1 port map( A1 => n200, A2 => n201, A3 => n202, ZN => n197);
   U478 : NAND3_X1 port map( A1 => n354, A2 => n455, A3 => n485, ZN => n353);
   U480 : NAND3_X1 port map( A1 => n554, A2 => n515, A3 => n633, ZN => n432);
   U483 : NAND3_X1 port map( A1 => r2(0), A2 => n469, A3 => r2(4), ZN => n86);
   U3 : INV_X1 port map( A => n667, ZN => n455);
   U4 : NAND3_X1 port map( A1 => n469, A2 => n672, A3 => r2(4), ZN => n168);
   U5 : AOI221_X1 port map( B1 => n637, B2 => r1(24), C1 => n638, C2 => r1(25),
                           A => n209, ZN => n208);
   U6 : NOR2_X1 port map( A1 => n671, A2 => r2(2), ZN => n437);
   U7 : AOI221_X1 port map( B1 => r1(22), B2 => n641, C1 => r1(23), C2 => n457,
                           A => n210, ZN => n207);
   U8 : AND2_X1 port map( A1 => n366, A2 => n530, ZN => n471);
   U9 : INV_X1 port map( A => n355, ZN => n653);
   U10 : NAND2_X1 port map( A1 => n669, A2 => n433, ZN => n355);
   U11 : INV_X1 port map( A => n286, ZN => n659);
   U12 : NAND3_X1 port map( A1 => n291, A2 => n161, A3 => n334, ZN => n160);
   U13 : BUF_X1 port map( A => n107, Z => n528);
   U14 : OAI221_X1 port map( B1 => n548, B2 => n674, C1 => n539, C2 => n675, A 
                           => n191, ZN => n189);
   U15 : OAI222_X1 port map( A1 => n673, A2 => n167, B1 => n168, B2 => n677, C1
                           => n676, C2 => n526, ZN => n190);
   U16 : NOR2_X1 port map( A1 => n670, A2 => r2(1), ZN => n442);
   U17 : OAI222_X1 port map( A1 => n676, A2 => n167, B1 => n168, B2 => n611, C1
                           => n619, C2 => n526, ZN => n166);
   U18 : AOI221_X1 port map( B1 => n604, B2 => n666, C1 => n601, C2 => n659, A 
                           => n147, ZN => n136);
   U19 : AOI221_X1 port map( B1 => n606, B2 => n666, C1 => n604, C2 => n659, A 
                           => n115, ZN => n96);
   U20 : INV_X1 port map( A => n471, ZN => n129);
   U21 : INV_X1 port map( A => n466, ZN => n363);
   U22 : AOI221_X1 port map( B1 => n592, B2 => n653, C1 => r1(6), C2 => n667, A
                           => n282, ZN => n275);
   U23 : AOI221_X1 port map( B1 => n586, B2 => n666, C1 => n581, C2 => n659, A 
                           => n240, ZN => n229);
   U24 : AOI221_X1 port map( B1 => n590, B2 => n666, C1 => n586, C2 => n659, A 
                           => n226, ZN => n215);
   U25 : AOI221_X1 port map( B1 => n592, B2 => n666, C1 => n590, C2 => n659, A 
                           => n203, ZN => n202);
   U26 : INV_X1 port map( A => n154, ZN => n664);
   U27 : OAI222_X1 port map( A1 => n569, A2 => n546, B1 => n431, B2 => n403, C1
                           => n576, C2 => n550, ZN => N1158);
   U28 : OAI221_X1 port map( B1 => n402, B2 => n403, C1 => n110, C2 => n557, A 
                           => n404, ZN => N1165);
   U29 : AOI221_X1 port map( B1 => n636, B2 => n560, C1 => n648, C2 => n557, A 
                           => n315, ZN => n381);
   U30 : AOI222_X1 port map( A1 => n648, A2 => n563, B1 => n359, B2 => n372, C1
                           => r1(2), C2 => n636, ZN => n371);
   U31 : BUF_X1 port map( A => n107, Z => n529);
   U32 : CLKBUF_X1 port map( A => n128, Z => n456);
   U33 : AND2_X1 port map( A1 => n351, A2 => n642, ZN => n457);
   U34 : OR3_X1 port map( A1 => r2(5), A2 => r2(31), A3 => r2(30), ZN => n458);
   U35 : AND2_X1 port map( A1 => n430, A2 => n471, ZN => n459);
   U36 : AND2_X1 port map( A1 => n103, A2 => n102, ZN => n460);
   U37 : OR3_X1 port map( A1 => r2(25), A2 => r2(24), A3 => r2(23), ZN => n461)
                           ;
   U38 : OR3_X1 port map( A1 => n188, A2 => n189, A3 => n190, ZN => n462);
   U39 : OR2_X1 port map( A1 => n518, A2 => n517, ZN => n463);
   U40 : OR2_X1 port map( A1 => n512, A2 => n511, ZN => n464);
   U41 : AND2_X1 port map( A1 => n111, A2 => n110, ZN => n364);
   U42 : AND4_X2 port map( A1 => n446, A2 => n467, A3 => n444, A4 => n445, ZN 
                           => n439);
   U43 : CLKBUF_X3 port map( A => n174, Z => n540);
   U44 : CLKBUF_X1 port map( A => n658, Z => n465);
   U45 : AND2_X1 port map( A1 => n113, A2 => n470, ZN => n390);
   U46 : BUF_X2 port map( A => n434, Z => n502);
   U47 : AND2_X2 port map( A1 => n439, A2 => n468, ZN => n434);
   U48 : NAND2_X1 port map( A1 => n196, A2 => n654, ZN => n315);
   U49 : INV_X1 port map( A => n86, ZN => n661);
   U50 : AND2_X2 port map( A1 => n437, A2 => n433, ZN => n466);
   U51 : NAND2_X1 port map( A1 => n661, A2 => n436, ZN => n116);
   U52 : NAND2_X1 port map( A1 => n661, A2 => n438, ZN => n100);
   U53 : NOR2_X1 port map( A1 => n448, A2 => n458, ZN => n467);
   U54 : AND2_X1 port map( A1 => n672, A2 => n668, ZN => n468);
   U55 : AND4_X2 port map( A1 => n447, A2 => n446, A3 => n444, A4 => n445, ZN 
                           => n469);
   U56 : AOI221_X1 port map( B1 => r1(22), B2 => n637, C1 => r1(23), C2 => n638
                           , A => n237, ZN => n236);
   U57 : NOR2_X1 port map( A1 => n187, A2 => n462, ZN => n185);
   U58 : NAND2_X1 port map( A1 => n502, A2 => n436, ZN => n366);
   U59 : OR2_X1 port map( A1 => n627, A2 => n494, ZN => n509);
   U60 : AND3_X1 port map( A1 => n283, A2 => n355, A3 => n168, ZN => n470);
   U61 : AND2_X1 port map( A1 => n524, A2 => n167, ZN => n443);
   U62 : INV_X1 port map( A => n167, ZN => n650);
   U63 : INV_X1 port map( A => n111, ZN => n652);
   U64 : NAND2_X1 port map( A1 => n632, A2 => n459, ZN => n429);
   U65 : NAND2_X1 port map( A1 => n666, A2 => r2(3), ZN => n472);
   U66 : AND3_X2 port map( A1 => n390, A2 => n364, A3 => n527, ZN => n351);
   U67 : NAND2_X2 port map( A1 => n435, A2 => n502, ZN => n110);
   U68 : AND3_X1 port map( A1 => n364, A2 => n390, A3 => n527, ZN => n473);
   U69 : AND3_X1 port map( A1 => n364, A2 => n390, A3 => n527, ZN => n500);
   U70 : OR2_X1 port map( A1 => n627, A2 => n544, ZN => n474);
   U71 : OR2_X1 port map( A1 => n628, A2 => n550, ZN => n475);
   U72 : NAND3_X1 port map( A1 => n474, A2 => n475, A3 => n130, ZN => N1185);
   U73 : CLKBUF_X1 port map( A => n640, Z => n476);
   U74 : INV_X1 port map( A => n528, ZN => n640);
   U75 : AND2_X1 port map( A1 => n551, A2 => n657, ZN => n477);
   U76 : AND2_X1 port map( A1 => n664, A2 => n561, ZN => n478);
   U77 : NOR3_X1 port map( A1 => n477, A2 => n478, A3 => n228, ZN => n227);
   U78 : NAND2_X1 port map( A1 => n654, A2 => n231, ZN => n479);
   U79 : NAND2_X1 port map( A1 => n590, A2 => n655, ZN => n480);
   U80 : INV_X1 port map( A => n232, ZN => n481);
   U81 : AND3_X1 port map( A1 => n479, A2 => n480, A3 => n481, ZN => n230);
   U82 : INV_X1 port map( A => n199, ZN => n657);
   U83 : OR2_X1 port map( A1 => n84, A2 => n464, ZN => n629);
   U84 : NAND2_X1 port map( A1 => r1(26), A2 => n641, ZN => n482);
   U85 : NAND2_X1 port map( A1 => r1(27), A2 => n457, ZN => n483);
   U86 : INV_X1 port map( A => n109, ZN => n484);
   U87 : AND3_X1 port map( A1 => n482, A2 => n483, A3 => n484, ZN => n104);
   U88 : CLKBUF_X1 port map( A => n634, Z => n485);
   U89 : CLKBUF_X1 port map( A => n93, Z => n486);
   U90 : OR2_X1 port map( A1 => n588, A2 => n546, ZN => n487);
   U91 : OR2_X1 port map( A1 => n591, A2 => n550, ZN => n488);
   U92 : NAND3_X1 port map( A1 => n487, A2 => n488, A3 => n123, ZN => n452);
   U93 : AOI221_X1 port map( B1 => r1(16), B2 => n641, C1 => r1(17), C2 => n457
                           , A => n298, ZN => n295);
   U94 : AOI221_X1 port map( B1 => r1(20), B2 => n641, C1 => n618, C2 => n457, 
                           A => n238, ZN => n235);
   U95 : AOI221_X1 port map( B1 => n617, B2 => n641, C1 => r1(22), C2 => n457, 
                           A => n224, ZN => n221);
   U96 : NOR3_X1 port map( A1 => r2(11), A2 => r2(12), A3 => r2(10), ZN => n489
                           );
   U97 : NOR2_X1 port map( A1 => n451, A2 => n490, ZN => n444);
   U98 : INV_X1 port map( A => n489, ZN => n490);
   U99 : AND2_X1 port map( A1 => n491, A2 => n522, ZN => n445);
   U100 : NOR4_X1 port map( A1 => r2(20), A2 => r2(19), A3 => r2(22), A4 => 
                           r2(21), ZN => n491);
   U101 : OR2_X1 port map( A1 => n623, A2 => n540, ZN => n492);
   U102 : OR2_X1 port map( A1 => n538, A2 => n624, ZN => n493);
   U103 : NAND3_X1 port map( A1 => n193, A2 => n493, A3 => n492, ZN => n187);
   U104 : BUF_X2 port map( A => n175, Z => n538);
   U105 : NAND2_X1 port map( A1 => n515, A2 => n351, ZN => n494);
   U106 : NOR2_X2 port map( A1 => n153, A2 => n89, ZN => n196);
   U107 : OR2_X1 port map( A1 => n676, A2 => n545, ZN => n495);
   U108 : OR2_X1 port map( A1 => n619, A2 => n550, ZN => n496);
   U109 : NAND3_X1 port map( A1 => n495, A2 => n496, A3 => n284, ZN => N1176);
   U110 : NAND2_X1 port map( A1 => n579, A2 => n656, ZN => n497);
   U111 : NAND2_X1 port map( A1 => n291, A2 => n292, ZN => n498);
   U112 : NAND2_X1 port map( A1 => n571, A2 => n663, ZN => n499);
   U113 : AND3_X1 port map( A1 => n497, A2 => n498, A3 => n499, ZN => n290);
   U114 : INV_X1 port map( A => n100, ZN => n656);
   U115 : AND2_X1 port map( A1 => n521, A2 => n520, ZN => n501);
   U116 : AND2_X1 port map( A1 => n519, A2 => n501, ZN => n97);
   U117 : NOR2_X1 port map( A1 => n95, A2 => n463, ZN => n92);
   U118 : INV_X1 port map( A => n110, ZN => n645);
   U119 : OAI221_X4 port map( B1 => n111, B2 => n577, C1 => n110, C2 => n585, A
                           => n373, ZN => n372);
   U120 : AND2_X1 port map( A1 => n586, A2 => n657, ZN => n503);
   U121 : AND2_X1 port map( A1 => n590, A2 => n664, ZN => n504);
   U122 : NOR3_X1 port map( A1 => n135, A2 => n504, A3 => n503, ZN => n133);
   U123 : AND2_X1 port map( A1 => r1(27), A2 => n637, ZN => n505);
   U124 : AND2_X1 port map( A1 => n638, A2 => r1(28), ZN => n506);
   U125 : NOR3_X1 port map( A1 => n505, A2 => n506, A3 => n144, ZN => n143);
   U126 : NAND2_X1 port map( A1 => n667, A2 => n436, ZN => n117);
   U127 : INV_X2 port map( A => n283, ZN => n507);
   U128 : NAND2_X1 port map( A1 => r1(28), A2 => n637, ZN => n508);
   U129 : INV_X1 port map( A => n106, ZN => n510);
   U130 : AND3_X1 port map( A1 => n508, A2 => n510, A3 => n509, ZN => n105);
   U131 : AND2_X1 port map( A1 => r1(30), A2 => n646, ZN => n511);
   U132 : AND2_X1 port map( A1 => r1(31), A2 => n523, ZN => n512);
   U133 : NOR2_X1 port map( A1 => n448, A2 => n458, ZN => n447);
   U134 : CLKBUF_X1 port map( A => n364, Z => n513);
   U135 : INV_X1 port map( A => n124, ZN => n514);
   U136 : NAND3_X1 port map( A1 => n105, A2 => n104, A3 => n460, ZN => n98);
   U137 : INV_X1 port map( A => n531, ZN => n649);
   U138 : OR4_X2 port map( A1 => r2(7), A2 => r2(6), A3 => r2(8), A4 => r2(9), 
                           ZN => n448);
   U139 : NAND2_X1 port map( A1 => n666, A2 => r2(3), ZN => n120);
   U140 : AND2_X1 port map( A1 => n437, A2 => r2(3), ZN => n435);
   U141 : AND4_X2 port map( A1 => n128, A2 => n471, A3 => n443, A4 => n417, ZN 
                           => n515);
   U142 : AND2_X1 port map( A1 => r2(0), A2 => n668, ZN => n516);
   U143 : AND2_X2 port map( A1 => n439, A2 => n516, ZN => n433);
   U144 : AND2_X1 port map( A1 => n590, A2 => n657, ZN => n517);
   U145 : AND2_X1 port map( A1 => n592, A2 => n664, ZN => n518);
   U146 : NAND2_X1 port map( A1 => n98, A2 => n654, ZN => n519);
   U147 : NAND2_X1 port map( A1 => n542, A2 => n655, ZN => n520);
   U148 : INV_X1 port map( A => n99, ZN => n521);
   U149 : NOR3_X1 port map( A1 => r2(17), A2 => r2(18), A3 => r2(16), ZN => 
                           n522);
   U150 : INV_X2 port map( A => n289, ZN => n666);
   U151 : INV_X2 port map( A => n367, ZN => n642);
   U152 : INV_X2 port map( A => n101, ZN => n663);
   U153 : NOR2_X2 port map( A1 => n670, A2 => n671, ZN => n436);
   U154 : CLKBUF_X1 port map( A => n114, Z => n547);
   U155 : CLKBUF_X1 port map( A => r1(0), Z => n555);
   U156 : CLKBUF_X1 port map( A => r1(0), Z => n556);
   U157 : NOR2_X1 port map( A1 => n449, A2 => n461, ZN => n446);
   U158 : INV_X1 port map( A => n160, ZN => n654);
   U159 : INV_X1 port map( A => n315, ZN => n634);
   U160 : INV_X1 port map( A => n161, ZN => n655);
   U161 : INV_X1 port map( A => n534, ZN => n639);
   U162 : NOR2_X1 port map( A1 => n663, A2 => n656, ZN => n291);
   U163 : INV_X1 port map( A => n196, ZN => n631);
   U164 : NAND2_X1 port map( A1 => n196, A2 => n334, ZN => n270);
   U165 : NOR2_X1 port map( A1 => n557, A2 => n550, ZN => N1155);
   U166 : INV_X1 port map( A => n366, ZN => n643);
   U167 : INV_X1 port map( A => n117, ZN => n662);
   U168 : INV_X1 port map( A => n426, ZN => n632);
   U169 : AND4_X1 port map( A1 => n117, A2 => n116, A3 => n289, A4 => n286, ZN 
                           => n334);
   U170 : INV_X1 port map( A => n121, ZN => n646);
   U171 : NAND2_X1 port map( A1 => n437, A2 => n661, ZN => n161);
   U172 : NAND2_X1 port map( A1 => n437, A2 => n667, ZN => n101);
   U173 : OAI22_X1 port map( A1 => n100, A2 => n614, B1 => n101, B2 => n611, ZN
                           => n99);
   U174 : AOI22_X1 port map( A1 => n573, A2 => n666, B1 => r1(2), B2 => n659, 
                           ZN => n258);
   U175 : AOI22_X1 port map( A1 => n581, A2 => n666, B1 => n573, B2 => n659, ZN
                           => n245);
   U176 : INV_X1 port map( A => n554, ZN => n557);
   U177 : AOI22_X1 port map( A1 => n580, A2 => n657, B1 => n553, B2 => n465, ZN
                           => n155);
   U178 : AOI22_X1 port map( A1 => n573, A2 => n657, B1 => n665, B2 => n565, ZN
                           => n181);
   U179 : AOI22_X1 port map( A1 => n573, A2 => n665, B1 => n660, B2 => n565, ZN
                           => n151);
   U180 : OAI22_X1 port map( A1 => n560, A2 => n550, B1 => n557, B2 => n543, ZN
                           => N1156);
   U181 : NAND2_X1 port map( A1 => n442, A2 => n667, ZN => n289);
   U182 : NAND2_X1 port map( A1 => n442, A2 => n661, ZN => n286);
   U183 : INV_X1 port map( A => n582, ZN => n585);
   U184 : NAND2_X1 port map( A1 => n442, A2 => n434, ZN => n367);
   U185 : INV_X1 port map( A => n119, ZN => n665);
   U186 : NAND2_X1 port map( A1 => n667, A2 => n669, ZN => n94);
   U187 : NAND2_X1 port map( A1 => n434, A2 => n669, ZN => n283);
   U188 : INV_X1 port map( A => n403, ZN => n633);
   U189 : CLKBUF_X1 port map( A => n172, Z => n532);
   U190 : BUF_X1 port map( A => n121, Z => n543);
   U191 : CLKBUF_X1 port map( A => n121, Z => n544);
   U192 : CLKBUF_X1 port map( A => n108, Z => n535);
   U193 : CLKBUF_X1 port map( A => n172, Z => n533);
   U194 : CLKBUF_X1 port map( A => n121, Z => n545);
   U195 : CLKBUF_X1 port map( A => n121, Z => n546);
   U196 : INV_X1 port map( A => n118, ZN => n660);
   U197 : INV_X1 port map( A => n564, ZN => n560);
   U198 : AOI211_X1 port map( C1 => n137, C2 => n136, A => n657, B => n664, ZN 
                           => n135);
   U199 : AOI22_X1 port map( A1 => n590, A2 => n652, B1 => n592, B2 => n645, ZN
                           => n342);
   U200 : AOI22_X1 port map( A1 => n592, A2 => n652, B1 => n597, B2 => n645, ZN
                           => n332);
   U201 : OAI222_X1 port map( A1 => n118, A2 => n578, B1 => n119, B2 => n585, 
                           C1 => n569, C2 => n472, ZN => n132);
   U202 : AOI221_X1 port map( B1 => n592, B2 => n507, C1 => r1(6), C2 => n653, 
                           A => n299, ZN => n294);
   U203 : AOI221_X1 port map( B1 => n606, B2 => n507, C1 => n604, C2 => n653, A
                           => n239, ZN => n234);
   U204 : INV_X1 port map( A => n613, ZN => n614);
   U205 : OAI221_X1 port map( B1 => n324, B2 => n270, C1 => n325, C2 => n315, A
                           => n326, ZN => N1173);
   U206 : AOI22_X1 port map( A1 => n646, A2 => r1(17), B1 => n523, B2 => r1(18)
                           , ZN => n326);
   U207 : AOI22_X1 port map( A1 => n552, A2 => n663, B1 => n656, B2 => n562, ZN
                           => n324);
   U208 : NOR4_X1 port map( A1 => n327, A2 => n328, A3 => n329, A4 => n330, ZN 
                           => n325);
   U209 : INV_X1 port map( A => n601, ZN => n603);
   U210 : AOI22_X1 port map( A1 => n515, A2 => n561, B1 => n553, B2 => n466, ZN
                           => n431);
   U211 : OAI221_X1 port map( B1 => n540, B2 => n619, C1 => n538, C2 => n620, A
                           => n254, ZN => n248);
   U212 : AOI22_X1 port map( A1 => r1(17), A2 => n639, B1 => r1(18), B2 => n640
                           , ZN => n254);
   U213 : OAI221_X1 port map( B1 => n540, B2 => n611, C1 => n538, C2 => n614, A
                           => n352, ZN => n345);
   U214 : AOI22_X1 port map( A1 => n600, A2 => n639, B1 => n604, B2 => n476, ZN
                           => n352);
   U215 : INV_X1 port map( A => n610, ZN => n611);
   U216 : OAI22_X1 port map( A1 => n116, A2 => n568, B1 => n117, B2 => n576, ZN
                           => n240);
   U217 : OAI22_X1 port map( A1 => n116, A2 => n575, B1 => n117, B2 => n585, ZN
                           => n226);
   U218 : OAI221_X1 port map( B1 => n268, B2 => n631, C1 => n269, C2 => n270, A
                           => n271, ZN => N1177);
   U219 : AOI22_X1 port map( A1 => n646, A2 => n617, B1 => n523, B2 => r1(22), 
                           ZN => n271);
   U220 : AOI222_X1 port map( A1 => n551, A2 => n662, B1 => n565, B2 => n666, 
                           C1 => n659, C2 => n563, ZN => n268);
   U221 : AOI221_X1 port map( B1 => n579, B2 => n663, C1 => n573, C2 => n655, A
                           => n272, ZN => n269);
   U222 : OAI221_X1 port map( B1 => n560, B2 => n545, C1 => n570, C2 => n550, A
                           => n432, ZN => N1157);
   U223 : OAI221_X1 port map( B1 => n575, B2 => n545, C1 => n585, C2 => n550, A
                           => n429, ZN => N1159);
   U224 : OAI221_X1 port map( B1 => n677, B2 => n544, C1 => n611, C2 => n550, A
                           => n379, ZN => N1168);
   U225 : NAND4_X1 port map( A1 => n355, A2 => n455, A3 => n380, A4 => n381, ZN
                           => n379);
   U226 : AOI21_X1 port map( B1 => n359, B2 => n382, A => n507, ZN => n380);
   U227 : OAI221_X1 port map( B1 => n611, B2 => n545, C1 => n614, C2 => n550, A
                           => n369, ZN => N1169);
   U228 : NAND4_X1 port map( A1 => n485, A2 => n370, A3 => n355, A4 => n455, ZN
                           => n369);
   U229 : OAI22_X1 port map( A1 => n283, A2 => n557, B1 => n507, B2 => n371, ZN
                           => n370);
   U230 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n543, ZN => n87);
   U231 : NAND2_X1 port map( A1 => n435, A2 => n661, ZN => n118);
   U232 : AOI22_X1 port map( A1 => n586, A2 => n663, B1 => r1(6), B2 => n656, 
                           ZN => n260);
   U233 : INV_X1 port map( A => n578, ZN => n573);
   U234 : INV_X1 port map( A => n568, ZN => n565);
   U235 : NAND2_X1 port map( A1 => n435, A2 => n667, ZN => n119);
   U236 : INV_X1 port map( A => n598, ZN => n599);
   U237 : NAND2_X1 port map( A1 => n440, A2 => n667, ZN => n154);
   U238 : AOI21_X1 port map( B1 => n636, B2 => n574, A => n507, ZN => n358);
   U239 : AOI22_X1 port map( A1 => r1(17), A2 => n652, B1 => r1(18), B2 => n645
                           , ZN => n192);
   U240 : NAND4_X1 port map( A1 => n120, A2 => n94, A3 => n118, A4 => n441, ZN 
                           => n93);
   U241 : NOR2_X1 port map( A1 => n665, A2 => n658, ZN => n441);
   U242 : AOI22_X1 port map( A1 => n581, A2 => n667, B1 => n606, B2 => n650, ZN
                           => n309);
   U243 : AOI22_X1 port map( A1 => n600, A2 => n507, B1 => n597, B2 => n653, ZN
                           => n265);
   U244 : AOI22_X1 port map( A1 => n590, A2 => n507, B1 => n586, B2 => n653, ZN
                           => n310);
   U245 : AOI22_X1 port map( A1 => n612, A2 => n507, B1 => n610, B2 => n653, ZN
                           => n191);
   U246 : AOI22_X1 port map( A1 => n565, A2 => n507, B1 => n653, B2 => n562, ZN
                           => n349);
   U247 : OAI211_X1 port map( C1 => n363, C2 => n585, A => n471, B => n424, ZN 
                           => n423);
   U248 : INV_X1 port map( A => r2(1), ZN => n671);
   U249 : AND2_X1 port map( A1 => n434, A2 => n438, ZN => n523);
   U250 : INV_X1 port map( A => r2(2), ZN => n670);
   U251 : INV_X1 port map( A => n85, ZN => n669);
   U252 : BUF_X1 port map( A => n556, Z => n551);
   U253 : BUF_X1 port map( A => n583, Z => n581);
   U254 : INV_X1 port map( A => n134, ZN => n658);
   U255 : NAND2_X1 port map( A1 => n440, A2 => n661, ZN => n199);
   U256 : BUF_X1 port map( A => n555, Z => n553);
   U257 : BUF_X1 port map( A => n584, Z => n580);
   U258 : BUF_X1 port map( A => n584, Z => n579);
   U259 : BUF_X1 port map( A => n556, Z => n552);
   U260 : BUF_X1 port map( A => n555, Z => n554);
   U261 : BUF_X1 port map( A => n583, Z => n582);
   U262 : AOI221_X1 port map( B1 => n592, B2 => n649, C1 => n596, C2 => n642, A
                           => n395, ZN => n391);
   U263 : OAI22_X1 port map( A1 => n528, A2 => n673, B1 => n535, B2 => n616, ZN
                           => n237);
   U264 : AOI22_X1 port map( A1 => n560, A2 => n651, B1 => n417, B2 => n418, ZN
                           => n416);
   U265 : INV_X1 port map( A => n605, ZN => n604);
   U266 : NOR3_X1 port map( A1 => r2(2), A2 => r2(3), A3 => r2(1), ZN => n438);
   U267 : INV_X1 port map( A => n587, ZN => n586);
   U268 : OAI221_X1 port map( B1 => n366, B2 => n603, C1 => n367, C2 => n607, A
                           => n368, ZN => n361);
   U269 : AOI22_X1 port map( A1 => n608, A2 => n652, B1 => n613, B2 => n645, ZN
                           => n253);
   U270 : AOI22_X1 port map( A1 => n600, A2 => n652, B1 => n604, B2 => n645, ZN
                           => n311);
   U271 : INV_X1 port map( A => n607, ZN => n606);
   U272 : AOI22_X1 port map( A1 => n586, A2 => n652, B1 => r1(6), B2 => n645, 
                           ZN => n350);
   U273 : AOI22_X1 port map( A1 => n596, A2 => n652, B1 => n602, B2 => n645, ZN
                           => n322);
   U274 : INV_X1 port map( A => n594, ZN => n592);
   U275 : NOR4_X1 port map( A1 => n261, A2 => n262, A3 => n263, A4 => n264, ZN 
                           => n259);
   U276 : OAI221_X1 port map( B1 => n547, B2 => n607, C1 => n539, C2 => n605, A
                           => n265, ZN => n263);
   U277 : NOR4_X1 port map( A1 => n163, A2 => n164, A3 => n165, A4 => n166, ZN 
                           => n159);
   U278 : OAI221_X1 port map( B1 => n547, B2 => n615, C1 => n539, C2 => n674, A
                           => n170, ZN => n165);
   U279 : OAI222_X1 port map( A1 => n585, A2 => n545, B1 => n425, B2 => n426, 
                           C1 => n588, C2 => n550, ZN => N1160);
   U280 : AOI22_X1 port map( A1 => n456, A2 => n574, B1 => n466, B2 => n567, ZN
                           => n428);
   U281 : OAI222_X1 port map( A1 => n605, A2 => n544, B1 => n396, B2 => n397, 
                           C1 => n607, C2 => n550, ZN => N1166);
   U282 : OAI22_X1 port map( A1 => n116, A2 => n599, B1 => n117, B2 => n603, ZN
                           => n115);
   U283 : OAI222_X1 port map( A1 => n675, A2 => n543, B1 => n344, B2 => n315, 
                           C1 => n674, C2 => n550, ZN => N1171);
   U284 : NOR4_X1 port map( A1 => n345, A2 => n346, A3 => n347, A4 => n348, ZN 
                           => n344);
   U285 : OAI221_X1 port map( B1 => n548, B2 => n585, C1 => n539, C2 => n577, A
                           => n349, ZN => n347);
   U286 : AOI221_X1 port map( B1 => n586, B2 => n651, C1 => r1(6), C2 => n643, 
                           A => n394, ZN => n392);
   U287 : AOI221_X1 port map( B1 => n656, B2 => n577, C1 => n663, C2 => n566, A
                           => n304, ZN => n303);
   U288 : NOR4_X1 port map( A1 => n305, A2 => n306, A3 => n307, A4 => n308, ZN 
                           => n304);
   U289 : OAI221_X1 port map( B1 => n114, B2 => n599, C1 => n539, C2 => n593, A
                           => n310, ZN => n307);
   U290 : AOI221_X1 port map( B1 => n542, B2 => n507, C1 => n606, C2 => n653, A
                           => n225, ZN => n220);
   U291 : INV_X1 port map( A => n591, ZN => n590);
   U292 : OAI222_X1 port map( A1 => n118, A2 => n585, B1 => n119, B2 => n589, 
                           C1 => n472, C2 => n574, ZN => n90);
   U293 : OAI221_X1 port map( B1 => n246, B2 => n160, C1 => n161, C2 => n588, A
                           => n247, ZN => n243);
   U294 : AOI22_X1 port map( A1 => n590, A2 => n663, B1 => n592, B2 => n656, ZN
                           => n247);
   U295 : NOR4_X1 port map( A1 => n248, A2 => n249, A3 => n250, A4 => n251, ZN 
                           => n246);
   U296 : OAI222_X1 port map( A1 => n675, A2 => n167, B1 => n455, B2 => n599, 
                           C1 => n674, C2 => n525, ZN => n251);
   U297 : OAI221_X1 port map( B1 => n540, B2 => n615, C1 => n538, C2 => n616, A
                           => n312, ZN => n305);
   U298 : AOI22_X1 port map( A1 => n608, A2 => n639, B1 => n613, B2 => n640, ZN
                           => n312);
   U299 : OAI221_X1 port map( B1 => n540, B2 => n624, C1 => n538, C2 => n625, A
                           => n176, ZN => n163);
   U300 : AOI22_X1 port map( A1 => r1(22), A2 => n639, B1 => r1(23), B2 => n640
                           , ZN => n176);
   U301 : OAI221_X1 port map( B1 => n540, B2 => n614, C1 => n538, C2 => n675, A
                           => n343, ZN => n337);
   U302 : AOI22_X1 port map( A1 => n604, A2 => n639, B1 => n606, B2 => n476, ZN
                           => n343);
   U303 : OAI221_X1 port map( B1 => n540, B2 => n675, C1 => n538, C2 => n674, A
                           => n333, ZN => n327);
   U304 : AOI22_X1 port map( A1 => n606, A2 => n639, B1 => n542, B2 => n476, ZN
                           => n333);
   U305 : OAI221_X1 port map( B1 => n540, B2 => n674, C1 => n538, C2 => n615, A
                           => n323, ZN => n317);
   U306 : AOI22_X1 port map( A1 => n542, A2 => n639, B1 => n609, B2 => n476, ZN
                           => n323);
   U307 : AOI22_X1 port map( A1 => n617, A2 => n639, B1 => r1(22), B2 => n640, 
                           ZN => n193);
   U308 : INV_X1 port map( A => n542, ZN => n677);
   U309 : OAI22_X1 port map( A1 => n116, A2 => n593, B1 => n117, B2 => n599, ZN
                           => n147);
   U310 : OAI22_X1 port map( A1 => n116, A2 => n585, B1 => n117, B2 => n587, ZN
                           => n203);
   U311 : OAI221_X1 port map( B1 => n366, B2 => n589, C1 => n367, C2 => n594, A
                           => n401, ZN => n398);
   U312 : OAI221_X1 port map( B1 => n366, B2 => n595, C1 => n367, C2 => n603, A
                           => n386, ZN => n383);
   U313 : OAI221_X1 port map( B1 => n673, B2 => n543, C1 => n676, C2 => n550, A
                           => n300, ZN => N1175);
   U314 : NAND4_X1 port map( A1 => n301, A2 => n286, A3 => n117, A4 => n116, ZN
                           => n300);
   U315 : AOI221_X1 port map( B1 => n302, B2 => n289, C1 => n666, C2 => n557, A
                           => n631, ZN => n301);
   U316 : OAI22_X1 port map( A1 => n564, A2 => n161, B1 => n655, B2 => n303, ZN
                           => n302);
   U317 : NAND4_X1 port map( A1 => n196, A2 => n285, A3 => n117, A4 => n116, ZN
                           => n284);
   U318 : OAI22_X1 port map( A1 => n286, A2 => n557, B1 => n287, B2 => n659, ZN
                           => n285);
   U319 : AOI22_X1 port map( A1 => n288, A2 => n289, B1 => n666, B2 => n562, ZN
                           => n287);
   U320 : OAI221_X1 port map( B1 => n607, B2 => n546, C1 => n677, C2 => n550, A
                           => n387, ZN => N1167);
   U321 : NOR2_X1 port map( A1 => n548, A2 => n557, ZN => n389);
   U322 : AOI221_X1 port map( B1 => n652, B2 => n560, C1 => n391, C2 => n392, A
                           => n393, ZN => n388);
   U323 : OAI221_X1 port map( B1 => n622, B2 => n544, C1 => n623, C2 => n550, A
                           => n227, ZN => N1180);
   U324 : AOI21_X1 port map( B1 => n229, B2 => n230, A => n631, ZN => n228);
   U325 : OAI221_X1 port map( B1 => n593, B2 => n544, C1 => n599, C2 => n550, A
                           => n414, ZN => N1163);
   U326 : INV_X1 port map( A => n416, ZN => n635);
   U327 : AOI22_X1 port map( A1 => n643, A2 => n557, B1 => n126, B2 => n127, ZN
                           => n125);
   U328 : AOI21_X1 port map( B1 => n573, B2 => n466, A => n129, ZN => n126);
   U329 : OAI221_X1 port map( B1 => n614, B2 => n543, C1 => n675, C2 => n550, A
                           => n353, ZN => N1170);
   U330 : OAI22_X1 port map( A1 => n355, A2 => n557, B1 => n653, B2 => n356, ZN
                           => n354);
   U331 : AOI22_X1 port map( A1 => n357, A2 => n358, B1 => n507, B2 => n562, ZN
                           => n356);
   U332 : OAI221_X1 port map( B1 => n591, B2 => n543, C1 => n595, C2 => n550, A
                           => n420, ZN => N1162);
   U333 : OAI211_X1 port map( C1 => n553, C2 => n417, A => n633, B => n421, ZN 
                           => n420);
   U334 : INV_X1 port map( A => n87, ZN => n647);
   U335 : INV_X1 port map( A => n89, ZN => n630);
   U336 : OAI221_X1 port map( B1 => n599, B2 => n546, C1 => n603, C2 => n550, A
                           => n409, ZN => N1164);
   U337 : OAI21_X1 port map( B1 => n410, B2 => n411, A => n633, ZN => n409);
   U338 : OAI221_X1 port map( B1 => n366, B2 => n574, C1 => n530, C2 => n585, A
                           => n412, ZN => n411);
   U339 : OAI221_X1 port map( B1 => n620, B2 => n546, C1 => n621, C2 => n550, A
                           => n255, ZN => N1178);
   U340 : OAI21_X1 port map( B1 => n256, B2 => n257, A => n196, ZN => n255);
   U341 : OAI221_X1 port map( B1 => n560, B2 => n117, C1 => n116, C2 => n557, A
                           => n258, ZN => n257);
   U342 : OAI221_X1 port map( B1 => n259, B2 => n160, C1 => n161, C2 => n585, A
                           => n260, ZN => n256);
   U343 : OAI22_X1 port map( A1 => n161, A2 => n568, B1 => n655, B2 => n290, ZN
                           => n288);
   U344 : NAND4_X1 port map( A1 => n293, A2 => n294, A3 => n295, A4 => n296, ZN
                           => n292);
   U345 : NOR3_X1 port map( A1 => n273, A2 => n663, A3 => n655, ZN => n272);
   U346 : OAI21_X1 port map( B1 => n586, B2 => n100, A => n274, ZN => n273);
   U347 : NAND4_X1 port map( A1 => n275, A2 => n276, A3 => n277, A4 => n278, ZN
                           => n274);
   U348 : OAI211_X1 port map( C1 => n624, C2 => n550, A => n212, B => n213, ZN 
                           => N1181);
   U350 : AOI22_X1 port map( A1 => n551, A2 => n665, B1 => n646, B2 => r1(25), 
                           ZN => n212);
   U351 : AOI221_X1 port map( B1 => n657, B2 => n563, C1 => n565, C2 => n664, A
                           => n214, ZN => n213);
   U352 : AOI21_X1 port map( B1 => n215, B2 => n216, A => n631, ZN => n214);
   U353 : OAI211_X1 port map( C1 => n625, C2 => n550, A => n194, B => n195, ZN 
                           => N1182);
   U354 : AOI22_X1 port map( A1 => n551, A2 => n660, B1 => n646, B2 => r1(26), 
                           ZN => n194);
   U355 : AOI221_X1 port map( B1 => n196, B2 => n197, C1 => n573, C2 => n664, A
                           => n198, ZN => n195);
   U356 : OAI22_X1 port map( A1 => n560, A2 => n119, B1 => n199, B2 => n569, ZN
                           => n198);
   U357 : AOI221_X1 port map( B1 => n138, B2 => n654, C1 => n606, C2 => n655, A
                           => n139, ZN => n137);
   U358 : OAI22_X1 port map( A1 => n611, A2 => n100, B1 => n677, B2 => n101, ZN
                           => n139);
   U359 : NAND2_X1 port map( A1 => r2(3), A2 => n436, ZN => n85);
   U360 : OAI22_X1 port map( A1 => n622, A2 => n529, B1 => n534, B2 => n621, ZN
                           => n144);
   U361 : AOI22_X1 port map( A1 => n604, A2 => n663, B1 => r1(11), B2 => n656, 
                           ZN => n186);
   U362 : AOI22_X1 port map( A1 => n606, A2 => n663, B1 => n656, B2 => n542, ZN
                           => n162);
   U363 : OAI22_X1 port map( A1 => n626, A2 => n550, B1 => n177, B2 => n89, ZN 
                           => N1183);
   U364 : AOI211_X1 port map( C1 => n646, C2 => r1(27), A => n179, B => n178, 
                           ZN => n177);
   U365 : OAI22_X1 port map( A1 => n472, A2 => n557, B1 => n560, B2 => n118, ZN
                           => n179);
   U366 : OAI221_X1 port map( B1 => n180, B2 => n153, C1 => n154, C2 => n585, A
                           => n181, ZN => n178);
   U368 : OAI22_X1 port map( A1 => n627, A2 => n550, B1 => n148, B2 => n89, ZN 
                           => N1184);
   U369 : NOR2_X1 port map( A1 => n149, A2 => n150, ZN => n148);
   U370 : OAI221_X1 port map( B1 => n560, B2 => n472, C1 => n626, C2 => n544, A
                           => n151, ZN => n150);
   U371 : OAI221_X1 port map( B1 => n152, B2 => n153, C1 => n154, C2 => n587, A
                           => n155, ZN => n149);
   U372 : AOI22_X1 port map( A1 => n542, A2 => n652, B1 => n609, B2 => n645, ZN
                           => n266);
   U373 : AND3_X1 port map( A1 => n671, A2 => n670, A3 => r2(3), ZN => n440);
   U374 : AOI221_X1 port map( B1 => n654, B2 => n217, C1 => n592, C2 => n655, A
                           => n218, ZN => n216);
   U375 : OAI22_X1 port map( A1 => n100, A2 => n603, B1 => n101, B2 => n599, ZN
                           => n218);
   U376 : NAND4_X1 port map( A1 => n219, A2 => n220, A3 => n221, A4 => n222, ZN
                           => n217);
   U377 : AOI222_X1 port map( A1 => n644, A2 => r1(18), B1 => n604, B2 => n667,
                           C1 => n650, C2 => r1(17), ZN => n219);
   U378 : NAND2_X1 port map( A1 => n659, A2 => r2(3), ZN => n134);
   U379 : NOR2_X1 port map( A1 => n182, A2 => n183, ZN => n180);
   U380 : OAI221_X1 port map( B1 => n117, B2 => n591, C1 => n116, C2 => n589, A
                           => n184, ZN => n183);
   U381 : OAI221_X1 port map( B1 => n185, B2 => n160, C1 => n161, C2 => n603, A
                           => n186, ZN => n182);
   U382 : AOI22_X1 port map( A1 => n596, A2 => n666, B1 => n592, B2 => n659, ZN
                           => n184);
   U383 : INV_X1 port map( A => r1(22), ZN => n620);
   U384 : NOR2_X1 port map( A1 => n156, A2 => n157, ZN => n152);
   U385 : OAI221_X1 port map( B1 => n117, B2 => n594, C1 => n116, C2 => n591, A
                           => n158, ZN => n157);
   U386 : OAI221_X1 port map( B1 => n159, B2 => n160, C1 => n161, C2 => n605, A
                           => n162, ZN => n156);
   U387 : AOI22_X1 port map( A1 => n601, A2 => n666, B1 => n597, B2 => n659, ZN
                           => n158);
   U388 : CLKBUF_X1 port map( A => r1(9), Z => n601);
   U389 : AOI22_X1 port map( A1 => n601, A2 => n663, B1 => n604, B2 => n656, ZN
                           => n200);
   U390 : AOI22_X1 port map( A1 => n654, A2 => n204, B1 => n598, B2 => n655, ZN
                           => n201);
   U391 : BUF_X1 port map( A => n558, Z => n562);
   U392 : CLKBUF_X1 port map( A => r1(9), Z => n600);
   U393 : INV_X1 port map( A => r1(18), ZN => n616);
   U394 : BUF_X1 port map( A => r1(13), Z => n608);
   U395 : BUF_X1 port map( A => n559, Z => n564);
   U396 : BUF_X1 port map( A => n559, Z => n563);
   U397 : CLKBUF_X1 port map( A => r1(8), Z => n597);
   U398 : BUF_X1 port map( A => r1(13), Z => n609);
   U399 : CLKBUF_X1 port map( A => r1(8), Z => n598);
   U400 : BUF_X1 port map( A => r1(21), Z => n617);
   U401 : CLKBUF_X1 port map( A => r1(8), Z => n596);
   U402 : BUF_X1 port map( A => n558, Z => n561);
   U403 : BUF_X1 port map( A => r1(14), Z => n612);
   U404 : BUF_X1 port map( A => r1(14), Z => n613);
   U405 : INV_X1 port map( A => r2(4), ZN => n668);
   U406 : CLKBUF_X1 port map( A => r1(9), Z => n602);
   U407 : BUF_X1 port map( A => r1(13), Z => n610);
   U408 : BUF_X1 port map( A => r1(21), Z => n618);
   U409 : CLKBUF_X1 port map( A => r1(4), Z => n583);
   U410 : CLKBUF_X1 port map( A => r1(4), Z => n584);
   U411 : OAI221_X1 port map( B1 => n547, B2 => n677, C1 => n539, C2 => n607, A
                           => n252, ZN => n250);
   U412 : AOI22_X1 port map( A1 => n604, A2 => n507, B1 => n602, B2 => n653, ZN
                           => n252);
   U413 : OAI221_X1 port map( B1 => n549, B2 => n588, C1 => n539, C2 => n585, A
                           => n341, ZN => n339);
   U414 : AOI22_X1 port map( A1 => n573, A2 => n507, B1 => n565, B2 => n653, ZN
                           => n341);
   U415 : OAI221_X1 port map( B1 => n547, B2 => n591, C1 => n539, C2 => n588, A
                           => n331, ZN => n329);
   U416 : AOI22_X1 port map( A1 => n580, A2 => n507, B1 => n573, B2 => n653, ZN
                           => n331);
   U417 : OAI221_X1 port map( B1 => n548, B2 => n595, C1 => n539, C2 => n591, A
                           => n321, ZN => n319);
   U418 : AOI22_X1 port map( A1 => n586, A2 => n507, B1 => n581, B2 => n653, ZN
                           => n321);
   U419 : AOI221_X1 port map( B1 => n641, B2 => r1(25), C1 => n457, C2 => 
                           r1(26), A => n145, ZN => n142);
   U420 : OAI221_X1 port map( B1 => n366, B2 => n599, C1 => n531, C2 => n603, A
                           => n376, ZN => n375);
   U421 : AOI22_X1 port map( A1 => n646, A2 => n600, B1 => n523, B2 => n604, ZN
                           => n404);
   U422 : NOR2_X1 port map( A1 => n405, A2 => n406, ZN => n402);
   U423 : OAI221_X1 port map( B1 => n366, B2 => n585, C1 => n531, C2 => n588, A
                           => n407, ZN => n406);
   U424 : OAI22_X1 port map( A1 => n529, A2 => n675, B1 => n535, B2 => n614, ZN
                           => n297);
   U425 : OAI22_X1 port map( A1 => n529, A2 => n676, B1 => n534, B2 => n673, ZN
                           => n223);
   U426 : INV_X1 port map( A => r1(15), ZN => n675);
   U427 : INV_X1 port map( A => r1(19), ZN => n673);
   U428 : AOI221_X1 port map( B1 => r1(16), B2 => n640, C1 => n609, C2 => n650,
                           A => n280, ZN => n277);
   U429 : OAI22_X1 port map( A1 => n534, A2 => n675, B1 => n532, B2 => n616, ZN
                           => n280);
   U430 : OAI221_X1 port map( B1 => n313, B2 => n270, C1 => n314, C2 => n315, A
                           => n316, ZN => N1174);
   U431 : AOI22_X1 port map( A1 => n646, A2 => r1(18), B1 => n523, B2 => r1(19)
                           , ZN => n316);
   U432 : AOI222_X1 port map( A1 => n565, A2 => n656, B1 => n552, B2 => n655, 
                           C1 => n663, C2 => n563, ZN => n313);
   U433 : NOR4_X1 port map( A1 => n317, A2 => n318, A3 => n319, A4 => n320, ZN 
                           => n314);
   U434 : AOI22_X1 port map( A1 => r1(18), A2 => n652, B1 => r1(19), B2 => n645
                           , ZN => n173);
   U435 : OAI221_X1 port map( B1 => n540, B2 => n676, C1 => n538, C2 => n619, A
                           => n267, ZN => n261);
   U436 : AOI22_X1 port map( A1 => r1(16), A2 => n639, B1 => r1(17), B2 => n640
                           , ZN => n267);
   U437 : INV_X1 port map( A => r1(20), ZN => n676);
   U438 : AOI221_X1 port map( B1 => r1(16), B2 => n507, C1 => r1(15), C2 => 
                           n653, A => n146, ZN => n141);
   U439 : INV_X1 port map( A => r1(16), ZN => n674);
   U440 : OAI221_X1 port map( B1 => n335, B2 => n315, C1 => n100, C2 => n557, A
                           => n336, ZN => N1172);
   U441 : AOI22_X1 port map( A1 => n646, A2 => r1(16), B1 => n523, B2 => r1(17)
                           , ZN => n336);
   U442 : NOR4_X1 port map( A1 => n337, A2 => n338, A3 => n339, A4 => n340, ZN 
                           => n335);
   U443 : OAI221_X1 port map( B1 => n241, B2 => n631, C1 => n154, C2 => n557, A
                           => n242, ZN => N1179);
   U444 : AOI22_X1 port map( A1 => n646, A2 => r1(23), B1 => n523, B2 => r1(24)
                           , ZN => n242);
   U445 : NOR2_X1 port map( A1 => n243, A2 => n244, ZN => n241);
   U446 : OAI221_X1 port map( B1 => n117, B2 => n567, C1 => n560, C2 => n116, A
                           => n245, ZN => n244);
   U447 : INV_X1 port map( A => r1(11), ZN => n607);
   U448 : OAI22_X1 port map( A1 => n528, A2 => n619, B1 => n535, B2 => n676, ZN
                           => n209);
   U449 : AOI22_X1 port map( A1 => r1(15), A2 => n507, B1 => n612, B2 => n653, 
                           ZN => n170);
   U450 : AOI221_X1 port map( B1 => r1(17), B2 => n507, C1 => r1(16), C2 => 
                           n653, A => n112, ZN => n103);
   U451 : NAND4_X1 port map( A1 => n205, A2 => n206, A3 => n207, A4 => n208, ZN
                           => n204);
   U452 : AOI222_X1 port map( A1 => n644, A2 => r1(19), B1 => n606, B2 => n667,
                           C1 => n650, C2 => r1(18), ZN => n205);
   U453 : AOI221_X1 port map( B1 => n608, B2 => n507, C1 => n542, C2 => n653, A
                           => n211, ZN => n206);
   U454 : OAI22_X1 port map( A1 => n100, A2 => n599, B1 => n101, B2 => n595, ZN
                           => n232);
   U455 : NAND4_X1 port map( A1 => n233, A2 => n234, A3 => n235, A4 => n236, ZN
                           => n231);
   U456 : AOI222_X1 port map( A1 => n644, A2 => r1(17), B1 => n601, B2 => n667,
                           C1 => n650, C2 => r1(16), ZN => n233);
   U457 : AOI221_X1 port map( B1 => r1(20), B2 => n638, C1 => r1(17), C2 => 
                           n641, A => n279, ZN => n278);
   U458 : OAI21_X1 port map( B1 => n540, B2 => n673, A => n100, ZN => n279);
   U459 : INV_X1 port map( A => r1(27), ZN => n625);
   U460 : INV_X1 port map( A => r1(28), ZN => n626);
   U461 : CLKBUF_X1 port map( A => r1(1), Z => n558);
   U462 : CLKBUF_X1 port map( A => r1(1), Z => n559);
   U463 : CLKBUF_X1 port map( A => r1(12), Z => n542);
   U464 : BUF_X1 port map( A => n113, Z => n539);
   U465 : INV_X1 port map( A => n113, ZN => n648);
   U466 : NAND2_X1 port map( A1 => n435, A2 => n433, ZN => n111);
   U467 : BUF_X1 port map( A => n169, Z => n524);
   U468 : CLKBUF_X1 port map( A => n169, Z => n525);
   U469 : CLKBUF_X1 port map( A => n169, Z => n526);
   U470 : NAND2_X1 port map( A1 => n440, A2 => n502, ZN => n169);
   U471 : OR3_X1 port map( A1 => r2(15), A2 => r2(14), A3 => r2(13), ZN => n451
                           );
   U472 : OAI22_X1 port map( A1 => n107, A2 => n623, B1 => n108, B2 => n622, ZN
                           => n106);
   U473 : INV_X1 port map( A => n494, ZN => n638);
   U474 : OAI221_X1 port map( B1 => n377, B2 => n677, C1 => n167, C2 => n587, A
                           => n378, ZN => n374);
   U475 : OAI221_X1 port map( B1 => n377, B2 => n599, C1 => n560, C2 => n167, A
                           => n408, ZN => n405);
   U479 : OAI221_X1 port map( B1 => n377, B2 => n595, C1 => n167, C2 => n557, A
                           => n413, ZN => n410);
   U481 : NAND4_X1 port map( A1 => n128, A2 => n471, A3 => n443, A4 => n417, ZN
                           => n377);
   U482 : OAI221_X1 port map( B1 => n398, B2 => n399, C1 => n564, C2 => n110, A
                           => n547, ZN => n396);
   U484 : OAI21_X1 port map( B1 => n565, B2 => n110, A => n549, ZN => n393);
   U485 : OAI222_X1 port map( A1 => n565, A2 => n111, B1 => n383, B2 => n384, 
                           C1 => n573, C2 => n110, ZN => n382);
   U486 : OAI222_X1 port map( A1 => n579, A2 => n111, B1 => n361, B2 => n362, 
                           C1 => n586, C2 => n110, ZN => n360);
   U487 : OAI22_X1 port map( A1 => n548, A2 => n605, B1 => n110, B2 => n677, ZN
                           => n281);
   U489 : OAI22_X1 port map( A1 => n110, A2 => n615, B1 => n111, B2 => n674, ZN
                           => n210);
   U490 : OAI22_X1 port map( A1 => n110, A2 => n674, B1 => n111, B2 => n675, ZN
                           => n224);
   U491 : OAI22_X1 port map( A1 => n110, A2 => n675, B1 => n111, B2 => n614, ZN
                           => n238);
   U492 : OAI22_X1 port map( A1 => n110, A2 => n607, B1 => n111, B2 => n605, ZN
                           => n298);
   U493 : OAI22_X1 port map( A1 => n676, A2 => n110, B1 => n111, B2 => n673, ZN
                           => n145);
   U494 : OAI22_X1 port map( A1 => n110, A2 => n619, B1 => n111, B2 => n676, ZN
                           => n109);
   U495 : NAND2_X1 port map( A1 => n642, A2 => r2(3), ZN => n527);
   U496 : BUF_X1 port map( A => n114, Z => n549);
   U497 : BUF_X1 port map( A => n114, Z => n548);
   U498 : INV_X1 port map( A => n114, ZN => n636);
   U499 : CLKBUF_X1 port map( A => n124, Z => n530);
   U500 : AOI221_X1 port map( B1 => r1(23), B2 => n637, C1 => n638, C2 => 
                           r1(24), A => n223, ZN => n222);
   U501 : AOI221_X1 port map( B1 => r1(18), B2 => n637, C1 => r1(19), C2 => 
                           n638, A => n297, ZN => n296);
   U502 : CLKBUF_X1 port map( A => n171, Z => n537);
   U503 : CLKBUF_X1 port map( A => n171, Z => n536);
   U504 : NAND2_X1 port map( A1 => n433, A2 => n438, ZN => n121);
   U505 : NAND2_X1 port map( A1 => n436, A2 => n433, ZN => n417);
   U506 : OAI211_X1 port map( C1 => n363, C2 => n677, A => n513, B => n365, ZN 
                           => n362);
   U507 : OAI21_X1 port map( B1 => n374, B2 => n375, A => n364, ZN => n373);
   U508 : OAI211_X1 port map( C1 => n363, C2 => n605, A => n513, B => n385, ZN 
                           => n384);
   U509 : OAI21_X1 port map( B1 => n363, B2 => n603, A => n513, ZN => n395);
   U510 : OAI211_X1 port map( C1 => n363, C2 => n599, A => n513, B => n400, ZN 
                           => n399);
   U511 : OAI211_X1 port map( C1 => n552, C2 => n525, A => n633, B => n415, ZN 
                           => n414);
   U512 : AOI21_X1 port map( B1 => n635, B2 => n526, A => n650, ZN => n415);
   U513 : NAND4_X1 port map( A1 => n633, A2 => n417, A3 => n167, A4 => n525, ZN
                           => n426);
   U514 : OAI222_X1 port map( A1 => n167, A2 => n603, B1 => n455, B2 => n570, 
                           C1 => n526, C2 => n605, ZN => n330);
   U515 : OAI222_X1 port map( A1 => n167, A2 => n605, B1 => n455, B2 => n578, 
                           C1 => n526, C2 => n607, ZN => n320);
   U516 : OAI222_X1 port map( A1 => n167, A2 => n599, B1 => n455, B2 => n560, 
                           C1 => n526, C2 => n603, ZN => n340);
   U517 : OAI222_X1 port map( A1 => n167, A2 => n595, B1 => n455, B2 => n557, 
                           C1 => n526, C2 => n599, ZN => n348);
   U518 : OAI222_X1 port map( A1 => n167, A2 => n577, B1 => n377, B2 => n605, 
                           C1 => n525, C2 => n585, ZN => n394);
   U519 : OAI222_X1 port map( A1 => n167, A2 => n614, B1 => n455, B2 => n595, 
                           C1 => n675, C2 => n525, ZN => n264);
   U520 : OAI211_X1 port map( C1 => n525, C2 => n677, A => n291, B => n309, ZN 
                           => n308);
   U521 : AOI22_X1 port map( A1 => n648, A2 => n566, B1 => n359, B2 => n360, ZN
                           => n357);
   U522 : NOR2_X1 port map( A1 => n636, A2 => n648, ZN => n359);
   U523 : NAND4_X1 port map( A1 => n143, A2 => n141, A3 => n142, A4 => n140, ZN
                           => n138);
   U524 : OAI211_X1 port map( C1 => n131, C2 => n132, A => n630, B => n647, ZN 
                           => n130);
   U525 : NAND2_X1 port map( A1 => n550, A2 => n469, ZN => n89);
   U526 : NAND2_X1 port map( A1 => n643, A2 => n473, ZN => n107);
   U527 : OAI222_X1 port map( A1 => n94, A2 => n557, B1 => n133, B2 => n486, C1
                           => n560, C2 => n134, ZN => n131);
   U528 : INV_X1 port map( A => n174, ZN => n637);
   U529 : AOI21_X1 port map( B1 => n642, B2 => n560, A => n129, ZN => n427);
   U530 : AOI222_X1 port map( A1 => n466, A2 => n560, B1 => n128, B2 => n567, 
                           C1 => n642, C2 => n557, ZN => n430);
   U531 : AOI22_X1 port map( A1 => n580, A2 => n456, B1 => r1(2), B2 => n642, 
                           ZN => n127);
   U532 : AOI22_X1 port map( A1 => n590, A2 => n642, B1 => n592, B2 => n466, ZN
                           => n407);
   U533 : AOI22_X1 port map( A1 => n586, A2 => n642, B1 => r1(6), B2 => n466, 
                           ZN => n412);
   U534 : AOI22_X1 port map( A1 => n573, A2 => n642, B1 => n586, B2 => n128, ZN
                           => n424);
   U535 : AOI222_X1 port map( A1 => n585, A2 => n642, B1 => n591, B2 => n128, 
                           C1 => n589, C2 => n466, ZN => n419);
   U536 : AOI22_X1 port map( A1 => n604, A2 => n642, B1 => n606, B2 => n466, ZN
                           => n376);
   U537 : NOR2_X1 port map( A1 => n466, A2 => n642, ZN => n128);
   U538 : NAND2_X1 port map( A1 => n642, A2 => r2(3), ZN => n114);
   U539 : CLKBUF_X1 port map( A => n124, Z => n531);
   U540 : NAND2_X1 port map( A1 => n442, A2 => n433, ZN => n124);
   U541 : NAND2_X1 port map( A1 => n634, A2 => n351, ZN => n403);
   U542 : NAND2_X1 port map( A1 => n351, A2 => n642, ZN => n172);
   U543 : BUF_X2 port map( A => n108, Z => n534);
   U544 : NAND2_X1 port map( A1 => n500, A2 => n651, ZN => n108);
   U545 : OR4_X2 port map( A1 => r2(27), A2 => r2(26), A3 => r2(29), A4 => 
                           r2(28), ZN => n449);
   U546 : NAND2_X1 port map( A1 => n515, A2 => n351, ZN => n175);
   U547 : AOI211_X1 port map( C1 => n422, C2 => n417, A => n644, B => n650, ZN 
                           => n421);
   U548 : AOI22_X1 port map( A1 => n565, A2 => n644, B1 => n573, B2 => n651, ZN
                           => n408);
   U549 : AOI22_X1 port map( A1 => n644, A2 => n561, B1 => r1(2), B2 => n651, 
                           ZN => n413);
   U550 : AOI222_X1 port map( A1 => n579, A2 => n651, B1 => n602, B2 => n515, 
                           C1 => n571, C2 => n644, ZN => n401);
   U551 : AOI221_X1 port map( B1 => n612, B2 => n644, C1 => n606, C2 => n652, A
                           => n281, ZN => n276);
   U552 : AOI222_X1 port map( A1 => n590, A2 => n651, B1 => n606, B2 => n515, 
                           C1 => r1(5), C2 => n644, ZN => n386);
   U553 : AOI222_X1 port map( A1 => n596, A2 => n651, B1 => n609, B2 => n515, 
                           C1 => r1(7), C2 => n644, ZN => n368);
   U554 : AOI22_X1 port map( A1 => n590, A2 => n644, B1 => n592, B2 => n651, ZN
                           => n378);
   U555 : AOI222_X1 port map( A1 => n608, A2 => n644, B1 => n586, B2 => n667, 
                           C1 => n542, C2 => n650, ZN => n293);
   U556 : AOI222_X1 port map( A1 => n644, A2 => r1(22), B1 => n612, B2 => n667,
                           C1 => n650, C2 => n617, ZN => n140);
   U557 : AOI222_X1 port map( A1 => r1(23), A2 => n644, B1 => r1(15), B2 => 
                           n667, C1 => r1(22), C2 => n650, ZN => n102);
   U558 : NAND2_X1 port map( A1 => n514, A2 => r2(3), ZN => n113);
   U559 : NAND2_X1 port map( A1 => n466, A2 => n351, ZN => n174);
   U560 : CLKBUF_X1 port map( A => n390, Z => n541);
   U561 : OAI22_X1 port map( A1 => n92, A2 => n486, B1 => n94, B2 => n560, ZN 
                           => n91);
   U562 : AOI211_X1 port map( C1 => n565, C2 => n465, A => n90, B => n91, ZN =>
                           n88);
   U563 : INV_X1 port map( A => r2(0), ZN => n672);
   U564 : AOI22_X1 port map( A1 => n427, A2 => n428, B1 => n553, B2 => n649, ZN
                           => n425);
   U565 : OAI211_X1 port map( C1 => n564, C2 => n530, A => n632, B => n125, ZN 
                           => n123);
   U566 : OAI221_X1 port map( B1 => n536, B2 => n611, C1 => n532, C2 => n614, A
                           => n332, ZN => n328);
   U567 : OAI221_X1 port map( B1 => n537, B2 => n614, C1 => n533, C2 => n675, A
                           => n322, ZN => n318);
   U568 : OAI221_X1 port map( B1 => n536, B2 => n677, C1 => n532, C2 => n611, A
                           => n342, ZN => n338);
   U569 : OAI221_X1 port map( B1 => n537, B2 => n607, C1 => n533, C2 => n677, A
                           => n350, ZN => n346);
   U570 : OAI221_X1 port map( B1 => n561, B2 => n366, C1 => n565, C2 => n531, A
                           => n423, ZN => n422);
   U571 : AOI22_X1 port map( A1 => n565, A2 => n650, B1 => r1(6), B2 => n649, 
                           ZN => n400);
   U572 : OAI221_X1 port map( B1 => n536, B2 => n673, C1 => n532, C2 => n676, A
                           => n253, ZN => n249);
   U573 : OAI222_X1 port map( A1 => n366, A2 => n565, B1 => n530, B2 => n573, 
                           C1 => n129, C2 => n419, ZN => n418);
   U574 : OAI221_X1 port map( B1 => n537, B2 => n616, C1 => n533, C2 => n673, A
                           => n266, ZN => n262);
   U575 : AOI22_X1 port map( A1 => n580, A2 => n650, B1 => n597, B2 => n649, ZN
                           => n385);
   U576 : OAI221_X1 port map( B1 => n622, B2 => n536, C1 => n623, C2 => n532, A
                           => n173, ZN => n164);
   U577 : AOI211_X1 port map( C1 => n97, C2 => n96, A => n657, B => n664, ZN =>
                           n95);
   U578 : OAI221_X1 port map( B1 => n537, B2 => n675, C1 => n533, C2 => n674, A
                           => n311, ZN => n306);
   U579 : AOI22_X1 port map( A1 => n590, A2 => n650, B1 => n604, B2 => n649, ZN
                           => n365);
   U580 : OAI221_X1 port map( B1 => n536, B2 => n621, C1 => n622, C2 => n533, A
                           => n192, ZN => n188);
   U581 : INV_X1 port map( A => n171, ZN => n641);
   U582 : NAND2_X1 port map( A1 => n473, A2 => n649, ZN => n171);
   U583 : OAI211_X1 port map( C1 => n552, C2 => n111, A => n541, B => n485, ZN 
                           => n397);
   U584 : OAI211_X1 port map( C1 => n388, C2 => n389, A => n541, B => n485, ZN 
                           => n387);
   U585 : OAI22_X1 port map( A1 => n283, A2 => n599, B1 => n539, B2 => n603, ZN
                           => n282);
   U586 : OAI22_X1 port map( A1 => n539, A2 => n614, B1 => n547, B2 => n675, ZN
                           => n211);
   U587 : OAI22_X1 port map( A1 => n539, A2 => n611, B1 => n547, B2 => n614, ZN
                           => n225);
   U588 : OAI22_X1 port map( A1 => n539, A2 => n677, B1 => n549, B2 => n611, ZN
                           => n239);
   U589 : OAI22_X1 port map( A1 => n539, A2 => n599, B1 => n114, B2 => n603, ZN
                           => n299);
   U590 : OAI22_X1 port map( A1 => n539, A2 => n615, B1 => n114, B2 => n616, ZN
                           => n146);
   U591 : OAI22_X1 port map( A1 => n539, A2 => n616, B1 => n114, B2 => n673, ZN
                           => n112);
   U592 : INV_X1 port map( A => n523, ZN => n550);
   U593 : INV_X1 port map( A => r1(2), ZN => n566);
   U594 : INV_X1 port map( A => r1(2), ZN => n567);
   U595 : INV_X1 port map( A => r1(2), ZN => n568);
   U596 : INV_X1 port map( A => r1(2), ZN => n569);
   U597 : INV_X1 port map( A => r1(2), ZN => n570);
   U598 : CLKBUF_X1 port map( A => r1(3), Z => n571);
   U599 : CLKBUF_X1 port map( A => r1(3), Z => n572);
   U600 : INV_X1 port map( A => n571, ZN => n574);
   U601 : INV_X1 port map( A => n571, ZN => n575);
   U602 : INV_X1 port map( A => n571, ZN => n576);
   U603 : INV_X1 port map( A => n572, ZN => n577);
   U604 : INV_X1 port map( A => r1(3), ZN => n578);
   U605 : INV_X1 port map( A => r1(5), ZN => n587);
   U606 : INV_X1 port map( A => r1(5), ZN => n588);
   U607 : INV_X1 port map( A => r1(5), ZN => n589);
   U608 : INV_X1 port map( A => r1(6), ZN => n591);
   U609 : INV_X1 port map( A => r1(7), ZN => n593);
   U610 : INV_X1 port map( A => r1(7), ZN => n594);
   U611 : INV_X1 port map( A => r1(7), ZN => n595);
   U612 : INV_X1 port map( A => r1(10), ZN => n605);
   U613 : INV_X1 port map( A => r1(17), ZN => n615);
   U614 : INV_X1 port map( A => n618, ZN => n619);
   U615 : INV_X1 port map( A => r1(23), ZN => n621);
   U616 : INV_X1 port map( A => r1(24), ZN => n622);
   U617 : INV_X1 port map( A => r1(25), ZN => n623);
   U618 : INV_X1 port map( A => r1(26), ZN => n624);
   U619 : INV_X1 port map( A => r1(29), ZN => n627);
   U620 : INV_X1 port map( A => r1(30), ZN => n628);
   U621 : INV_X2 port map( A => n524, ZN => n644);
   U622 : INV_X2 port map( A => n417, ZN => n651);
   U623 : INV_X2 port map( A => n168, ZN => n667);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity xor_gate_nbit32 is

   port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
         (31 downto 0));

end xor_gate_nbit32;

architecture SYN_beh of xor_gate_nbit32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B(9), B => A(9), Z => Y(9));
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => Y(8));
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => Y(7));
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => Y(6));
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => Y(5));
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => Y(4));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => Y(3));
   U8 : XOR2_X1 port map( A => B(31), B => A(31), Z => Y(31));
   U9 : XOR2_X1 port map( A => B(30), B => A(30), Z => Y(30));
   U10 : XOR2_X1 port map( A => B(2), B => A(2), Z => Y(2));
   U11 : XOR2_X1 port map( A => B(29), B => A(29), Z => Y(29));
   U12 : XOR2_X1 port map( A => B(28), B => A(28), Z => Y(28));
   U13 : XOR2_X1 port map( A => B(27), B => A(27), Z => Y(27));
   U14 : XOR2_X1 port map( A => B(26), B => A(26), Z => Y(26));
   U15 : XOR2_X1 port map( A => B(25), B => A(25), Z => Y(25));
   U16 : XOR2_X1 port map( A => B(24), B => A(24), Z => Y(24));
   U17 : XOR2_X1 port map( A => B(23), B => A(23), Z => Y(23));
   U18 : XOR2_X1 port map( A => B(22), B => A(22), Z => Y(22));
   U19 : XOR2_X1 port map( A => B(21), B => A(21), Z => Y(21));
   U20 : XOR2_X1 port map( A => B(20), B => A(20), Z => Y(20));
   U21 : XOR2_X1 port map( A => B(1), B => A(1), Z => Y(1));
   U22 : XOR2_X1 port map( A => B(19), B => A(19), Z => Y(19));
   U23 : XOR2_X1 port map( A => B(18), B => A(18), Z => Y(18));
   U24 : XOR2_X1 port map( A => B(17), B => A(17), Z => Y(17));
   U25 : XOR2_X1 port map( A => B(16), B => A(16), Z => Y(16));
   U26 : XOR2_X1 port map( A => B(15), B => A(15), Z => Y(15));
   U27 : XOR2_X1 port map( A => B(14), B => A(14), Z => Y(14));
   U28 : XOR2_X1 port map( A => B(13), B => A(13), Z => Y(13));
   U29 : XOR2_X1 port map( A => B(12), B => A(12), Z => Y(12));
   U30 : XOR2_X1 port map( A => B(11), B => A(11), Z => Y(11));
   U31 : XOR2_X1 port map( A => B(10), B => A(10), Z => Y(10));
   U32 : XOR2_X1 port map( A => B(0), B => A(0), Z => Y(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity or_gate_nbit32 is

   port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
         (31 downto 0));

end or_gate_nbit32;

architecture SYN_beh of or_gate_nbit32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A(31), A2 => B(31), ZN => Y(31));
   U2 : OR2_X1 port map( A1 => A(6), A2 => B(6), ZN => Y(6));
   U3 : OR2_X1 port map( A1 => A(4), A2 => B(4), ZN => Y(4));
   U4 : OR2_X1 port map( A1 => A(7), A2 => B(7), ZN => Y(7));
   U5 : OR2_X1 port map( A1 => A(9), A2 => B(9), ZN => Y(9));
   U6 : OR2_X1 port map( A1 => A(5), A2 => B(5), ZN => Y(5));
   U7 : OR2_X1 port map( A1 => A(3), A2 => B(3), ZN => Y(3));
   U8 : OR2_X1 port map( A1 => A(30), A2 => B(30), ZN => Y(30));
   U9 : OR2_X1 port map( A1 => A(21), A2 => B(21), ZN => Y(21));
   U10 : OR2_X1 port map( A1 => A(20), A2 => B(20), ZN => Y(20));
   U11 : OR2_X1 port map( A1 => A(29), A2 => B(29), ZN => Y(29));
   U12 : OR2_X1 port map( A1 => A(25), A2 => B(25), ZN => Y(25));
   U13 : OR2_X1 port map( A1 => A(26), A2 => B(26), ZN => Y(26));
   U14 : OR2_X1 port map( A1 => A(27), A2 => B(27), ZN => Y(27));
   U15 : OR2_X1 port map( A1 => A(23), A2 => B(23), ZN => Y(23));
   U16 : OR2_X1 port map( A1 => A(24), A2 => B(24), ZN => Y(24));
   U17 : OR2_X1 port map( A1 => A(15), A2 => B(15), ZN => Y(15));
   U18 : OR2_X1 port map( A1 => A(10), A2 => B(10), ZN => Y(10));
   U19 : OR2_X1 port map( A1 => A(13), A2 => B(13), ZN => Y(13));
   U20 : OR2_X1 port map( A1 => A(14), A2 => B(14), ZN => Y(14));
   U21 : OR2_X1 port map( A1 => A(11), A2 => B(11), ZN => Y(11));
   U22 : OR2_X1 port map( A1 => A(16), A2 => B(16), ZN => Y(16));
   U23 : OR2_X1 port map( A1 => A(12), A2 => B(12), ZN => Y(12));
   U24 : OR2_X1 port map( A1 => A(17), A2 => B(17), ZN => Y(17));
   U25 : OR2_X1 port map( A1 => A(18), A2 => B(18), ZN => Y(18));
   U26 : OR2_X1 port map( A1 => A(19), A2 => B(19), ZN => Y(19));
   U27 : OR2_X1 port map( A1 => A(1), A2 => B(1), ZN => Y(1));
   U28 : OR2_X1 port map( A1 => A(2), A2 => B(2), ZN => Y(2));
   U29 : OR2_X1 port map( A1 => A(22), A2 => B(22), ZN => Y(22));
   U30 : OR2_X1 port map( A1 => A(28), A2 => B(28), ZN => Y(28));
   U31 : OR2_X1 port map( A1 => A(0), A2 => B(0), ZN => Y(0));
   U32 : OR2_X1 port map( A1 => A(8), A2 => B(8), ZN => Y(8));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity and_gate_nbit32 is

   port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
         (31 downto 0));

end and_gate_nbit32;

architecture SYN_beh of and_gate_nbit32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => Y(5));
   U2 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => Y(12));
   U3 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => Y(7));
   U4 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => Y(9));
   U5 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => Y(6));
   U6 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => Y(4));
   U7 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => Y(3));
   U8 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => Y(31));
   U9 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => Y(17));
   U10 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => Y(14));
   U11 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => Y(23));
   U12 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => Y(11));
   U13 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => Y(18));
   U14 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => Y(1));
   U15 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => Y(15));
   U16 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => Y(27));
   U17 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => Y(16));
   U18 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => Y(24));
   U19 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => Y(21));
   U20 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => Y(10));
   U21 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => Y(25));
   U22 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => Y(19));
   U23 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => Y(20));
   U24 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => Y(13));
   U25 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => Y(26));
   U26 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => Y(29));
   U27 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => Y(30));
   U28 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => Y(2));
   U29 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => Y(22));
   U30 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => Y(28));
   U31 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => Y(0));
   U32 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => Y(8));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity P4_ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic;  Y : out std_logic_vector (31 downto 0));

end P4_ADDER_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32_NBIT_PER_BLOCK4_1 is

   component SUMGEN_NBIT32_NBLOCKS8_1
      port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
            std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal outCarryGen_7_port, outCarryGen_6_port, outCarryGen_5_port, 
      outCarryGen_4_port, outCarryGen_3_port, outCarryGen_2_port, 
      outCarryGen_1_port, outCarryGen_0_port : std_logic;

begin
   
   CG : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Cin => Cin, Co(7) 
                           => outCarryGen_7_port, Co(6) => outCarryGen_6_port, 
                           Co(5) => outCarryGen_5_port, Co(4) => 
                           outCarryGen_4_port, Co(3) => outCarryGen_3_port, 
                           Co(2) => outCarryGen_2_port, Co(1) => 
                           outCarryGen_1_port, Co(0) => outCarryGen_0_port);
   SG : SUMGEN_NBIT32_NBLOCKS8_1 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), cin_vect(7) => 
                           outCarryGen_7_port, cin_vect(6) => 
                           outCarryGen_6_port, cin_vect(5) => 
                           outCarryGen_5_port, cin_vect(4) => 
                           outCarryGen_4_port, cin_vect(3) => 
                           outCarryGen_3_port, cin_vect(2) => 
                           outCarryGen_2_port, cin_vect(1) => 
                           outCarryGen_1_port, cin_vect(0) => 
                           outCarryGen_0_port, Co => Cout, SUM(31) => Y(31), 
                           SUM(30) => Y(30), SUM(29) => Y(29), SUM(28) => Y(28)
                           , SUM(27) => Y(27), SUM(26) => Y(26), SUM(25) => 
                           Y(25), SUM(24) => Y(24), SUM(23) => Y(23), SUM(22) 
                           => Y(22), SUM(21) => Y(21), SUM(20) => Y(20), 
                           SUM(19) => Y(19), SUM(18) => Y(18), SUM(17) => Y(17)
                           , SUM(16) => Y(16), SUM(15) => Y(15), SUM(14) => 
                           Y(14), SUM(13) => Y(13), SUM(12) => Y(12), SUM(11) 
                           => Y(11), SUM(10) => Y(10), SUM(9) => Y(9), SUM(8) 
                           => Y(8), SUM(7) => Y(7), SUM(6) => Y(6), SUM(5) => 
                           Y(5), SUM(4) => Y(4), SUM(3) => Y(3), SUM(2) => Y(2)
                           , SUM(1) => Y(1), SUM(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n33, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n111, ZN => Y(0));
   U2 : INV_X1 port map( A => n122, ZN => Y(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n68, B1 => B(1), B2 => n74, ZN => 
                           n122);
   U4 : INV_X1 port map( A => n141, ZN => Y(8));
   U5 : INV_X1 port map( A => n142, ZN => Y(9));
   U6 : AOI22_X1 port map( A1 => A(9), A2 => n68, B1 => n77, B2 => B(9), ZN => 
                           n142);
   U7 : INV_X1 port map( A => n139, ZN => Y(6));
   U8 : AOI22_X1 port map( A1 => A(6), A2 => n69, B1 => B(6), B2 => n70, ZN => 
                           n139);
   U9 : INV_X1 port map( A => n124, ZN => Y(21));
   U10 : INV_X1 port map( A => n133, ZN => Y(2));
   U11 : AOI22_X1 port map( A1 => A(2), A2 => n69, B1 => B(2), B2 => n71, ZN =>
                           n133);
   U12 : INV_X1 port map( A => n121, ZN => Y(19));
   U13 : AOI22_X1 port map( A1 => A(19), A2 => n68, B1 => B(19), B2 => n75, ZN 
                           => n121);
   U14 : INV_X1 port map( A => n132, ZN => Y(29));
   U15 : AOI22_X1 port map( A1 => A(29), A2 => n69, B1 => B(29), B2 => n72, ZN 
                           => n132);
   U16 : INV_X1 port map( A => n78, ZN => n68);
   U17 : INV_X1 port map( A => n78, ZN => n69);
   U18 : INV_X1 port map( A => n112, ZN => Y(10));
   U19 : AOI22_X1 port map( A1 => A(10), A2 => n68, B1 => B(10), B2 => n77, ZN 
                           => n112);
   U20 : INV_X1 port map( A => n136, ZN => Y(3));
   U21 : AOI22_X1 port map( A1 => A(3), A2 => n68, B1 => B(3), B2 => n71, ZN =>
                           n136);
   U22 : INV_X1 port map( A => n129, ZN => Y(26));
   U23 : AOI22_X1 port map( A1 => A(26), A2 => n69, B1 => B(26), B2 => n72, ZN 
                           => n129);
   U24 : INV_X1 port map( A => n131, ZN => Y(28));
   U25 : INV_X1 port map( A => n137, ZN => Y(4));
   U26 : AOI22_X1 port map( A1 => A(4), A2 => n69, B1 => B(4), B2 => n71, ZN =>
                           n137);
   U27 : INV_X1 port map( A => n135, ZN => Y(31));
   U28 : AOI22_X1 port map( A1 => A(31), A2 => n68, B1 => B(31), B2 => n71, ZN 
                           => n135);
   U29 : INV_X1 port map( A => n113, ZN => Y(11));
   U30 : AOI22_X1 port map( A1 => A(11), A2 => n68, B1 => B(11), B2 => n77, ZN 
                           => n113);
   U31 : INV_X1 port map( A => n114, ZN => Y(12));
   U32 : AOI22_X1 port map( A1 => A(12), A2 => n68, B1 => B(12), B2 => n76, ZN 
                           => n114);
   U33 : INV_X1 port map( A => n115, ZN => Y(13));
   U34 : INV_X1 port map( A => n116, ZN => Y(14));
   U35 : AOI22_X1 port map( A1 => A(14), A2 => n68, B1 => B(14), B2 => n76, ZN 
                           => n116);
   U36 : INV_X1 port map( A => n117, ZN => Y(15));
   U37 : AOI22_X1 port map( A1 => A(15), A2 => n68, B1 => B(15), B2 => n76, ZN 
                           => n117);
   U38 : INV_X1 port map( A => n126, ZN => Y(23));
   U39 : AOI22_X1 port map( A1 => A(23), A2 => n69, B1 => B(23), B2 => n73, ZN 
                           => n126);
   U40 : INV_X1 port map( A => n119, ZN => Y(17));
   U41 : AOI22_X1 port map( A1 => A(17), A2 => n68, B1 => B(17), B2 => n75, ZN 
                           => n119);
   U42 : INV_X1 port map( A => n125, ZN => Y(22));
   U43 : INV_X1 port map( A => n118, ZN => Y(16));
   U44 : AOI22_X1 port map( A1 => A(16), A2 => n68, B1 => B(16), B2 => n75, ZN 
                           => n118);
   U45 : INV_X1 port map( A => n120, ZN => Y(18));
   U46 : AOI22_X1 port map( A1 => A(18), A2 => n68, B1 => B(18), B2 => n75, ZN 
                           => n120);
   U47 : INV_X1 port map( A => n138, ZN => Y(5));
   U48 : AOI22_X1 port map( A1 => A(5), A2 => n69, B1 => B(5), B2 => n70, ZN =>
                           n138);
   U49 : INV_X1 port map( A => n134, ZN => Y(30));
   U50 : AOI22_X1 port map( A1 => A(30), A2 => n69, B1 => B(30), B2 => n74, ZN 
                           => n134);
   U51 : INV_X1 port map( A => n130, ZN => Y(27));
   U52 : AOI22_X1 port map( A1 => A(27), A2 => n69, B1 => B(27), B2 => n72, ZN 
                           => n130);
   U53 : INV_X1 port map( A => n128, ZN => Y(25));
   U54 : AOI22_X1 port map( A1 => A(25), A2 => n69, B1 => B(25), B2 => n73, ZN 
                           => n128);
   U55 : INV_X1 port map( A => n123, ZN => Y(20));
   U56 : AOI22_X1 port map( A1 => A(20), A2 => n69, B1 => B(20), B2 => n74, ZN 
                           => n123);
   U57 : INV_X1 port map( A => n140, ZN => Y(7));
   U58 : AOI22_X1 port map( A1 => A(7), A2 => n68, B1 => B(7), B2 => n70, ZN =>
                           n140);
   U59 : INV_X1 port map( A => n127, ZN => Y(24));
   U60 : AOI22_X1 port map( A1 => A(24), A2 => n69, B1 => B(24), B2 => n73, ZN 
                           => n127);
   U61 : BUF_X1 port map( A => n66, Z => n75);
   U62 : BUF_X1 port map( A => n33, Z => n71);
   U63 : BUF_X1 port map( A => n67, Z => n78);
   U64 : BUF_X1 port map( A => n33, Z => n70);
   U65 : BUF_X1 port map( A => n67, Z => n76);
   U66 : BUF_X1 port map( A => n66, Z => n74);
   U67 : BUF_X1 port map( A => n33, Z => n72);
   U68 : BUF_X1 port map( A => n66, Z => n73);
   U69 : BUF_X1 port map( A => n67, Z => n77);
   U70 : BUF_X1 port map( A => SEL, Z => n66);
   U71 : BUF_X1 port map( A => SEL, Z => n67);
   U72 : BUF_X1 port map( A => SEL, Z => n33);
   U73 : AOI22_X1 port map( A1 => A(13), A2 => n68, B1 => B(13), B2 => n76, ZN 
                           => n115);
   U74 : AOI22_X1 port map( A1 => A(22), A2 => n69, B1 => B(22), B2 => n73, ZN 
                           => n125);
   U75 : AOI22_X1 port map( A1 => A(28), A2 => n69, B1 => B(28), B2 => n72, ZN 
                           => n131);
   U76 : AOI22_X1 port map( A1 => A(21), A2 => n69, B1 => B(21), B2 => n74, ZN 
                           => n124);
   U77 : AOI22_X1 port map( A1 => A(0), A2 => n68, B1 => B(0), B2 => n77, ZN =>
                           n111);
   U78 : AOI22_X1 port map( A1 => A(8), A2 => n69, B1 => B(8), B2 => n70, ZN =>
                           n141);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity SUMGEN_NBIT32_NBLOCKS8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
         std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
         std_logic_vector (31 downto 0));

end SUMGEN_NBIT32_NBLOCKS8_0;

architecture SYN_STRUCTURAL of SUMGEN_NBIT32_NBLOCKS8_0 is

   component CSblock_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component CSblock_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  cin : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133 : std_logic;

begin
   
   block_i_0 : CSblock_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), cin => cin_vect(0), Y(3) => 
                           SUM(3), Y(2) => SUM(2), Y(1) => SUM(1), Y(0) => 
                           SUM(0), Co => n_1127);
   block_i_1 : CSblock_NBIT4_31 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), cin => cin_vect(1), Y(3) => 
                           SUM(7), Y(2) => SUM(6), Y(1) => SUM(5), Y(0) => 
                           SUM(4), Co => n_1128);
   block_i_2 : CSblock_NBIT4_30 port map( A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), cin => cin_vect(2), Y(3)
                           => SUM(11), Y(2) => SUM(10), Y(1) => SUM(9), Y(0) =>
                           SUM(8), Co => n_1129);
   block_i_3 : CSblock_NBIT4_29 port map( A(3) => A(15), A(2) => A(14), A(1) =>
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), cin => cin_vect(3), 
                           Y(3) => SUM(15), Y(2) => SUM(14), Y(1) => SUM(13), 
                           Y(0) => SUM(12), Co => n_1130);
   block_i_4 : CSblock_NBIT4_28 port map( A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), cin => cin_vect(4), 
                           Y(3) => SUM(19), Y(2) => SUM(18), Y(1) => SUM(17), 
                           Y(0) => SUM(16), Co => n_1131);
   block_i_5 : CSblock_NBIT4_27 port map( A(3) => A(23), A(2) => A(22), A(1) =>
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), cin => cin_vect(5), 
                           Y(3) => SUM(23), Y(2) => SUM(22), Y(1) => SUM(21), 
                           Y(0) => SUM(20), Co => n_1132);
   block_i_6 : CSblock_NBIT4_26 port map( A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), cin => cin_vect(6), 
                           Y(3) => SUM(27), Y(2) => SUM(26), Y(1) => SUM(25), 
                           Y(0) => SUM(24), Co => n_1133);
   block_i_7 : CSblock_NBIT4_25 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), cin => cin_vect(7), 
                           Y(3) => SUM(31), Y(2) => SUM(30), Y(1) => SUM(29), 
                           Y(0) => SUM(28), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   component GENERAL_G_31
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_32
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_33
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_34
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_82
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_83
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_84
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_85
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_35
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_G_36
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_86
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_37
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_87
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_88
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_89
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_90
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_91
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_92
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_93
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_94
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_95
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_96
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_97
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_98
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_99
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_100
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_101
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_102
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_103
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_104
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_105
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_106
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_PG_107
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_38
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component GENERAL_PG_0
      port( G_in, P_in, G_in_prev, P_in_prev : in std_logic;  G_out, P_out : 
            out std_logic);
   end component;
   
   component GENERAL_G_39
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_97
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_98
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_99
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_100
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_101
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_102
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_103
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_104
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_105
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_106
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_107
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_108
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_109
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_110
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_111
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_112
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_113
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_114
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_115
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_116
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_117
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_118
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_119
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_120
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_121
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_122
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_123
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_124
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_125
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_126
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component PG_block_127
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   component GENERAL_G_0
      port( G_in, P_in, G_in_prev : in std_logic;  G_out : out std_logic);
   end component;
   
   component PG_block_0
      port( A, B : in std_logic;  G, P : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, first_generate, p_vett_4_3_port, p_vett_4_2_port, 
      p_vett_3_3_port, p_vett_3_2_port, p_vett_3_1_port, p_vett_2_7_port, 
      p_vett_2_6_port, p_vett_2_5_port, p_vett_2_4_port, p_vett_2_3_port, 
      p_vett_2_2_port, p_vett_2_1_port, p_vett_1_15_port, p_vett_1_14_port, 
      p_vett_1_13_port, p_vett_1_12_port, p_vett_1_11_port, p_vett_1_10_port, 
      p_vett_1_9_port, p_vett_1_8_port, p_vett_1_7_port, p_vett_1_6_port, 
      p_vett_1_5_port, p_vett_1_4_port, p_vett_1_3_port, p_vett_1_2_port, 
      p_vett_1_1_port, p_vett_0_31_port, p_vett_0_30_port, p_vett_0_29_port, 
      p_vett_0_28_port, p_vett_0_27_port, p_vett_0_26_port, p_vett_0_25_port, 
      p_vett_0_24_port, p_vett_0_23_port, p_vett_0_22_port, p_vett_0_21_port, 
      p_vett_0_20_port, p_vett_0_19_port, p_vett_0_18_port, p_vett_0_17_port, 
      p_vett_0_16_port, p_vett_0_15_port, p_vett_0_14_port, p_vett_0_13_port, 
      p_vett_0_12_port, p_vett_0_11_port, p_vett_0_10_port, p_vett_0_9_port, 
      p_vett_0_8_port, p_vett_0_7_port, p_vett_0_6_port, p_vett_0_5_port, 
      p_vett_0_4_port, p_vett_0_3_port, p_vett_0_2_port, p_vett_0_1_port, 
      p_vett_0_0_port, g_vett_4_3_port, g_vett_4_2_port, g_vett_3_3_port, 
      g_vett_3_2_port, g_vett_3_1_port, g_vett_2_7_port, g_vett_2_6_port, 
      g_vett_2_5_port, g_vett_2_4_port, g_vett_2_3_port, g_vett_2_2_port, 
      g_vett_2_1_port, g_vett_1_15_port, g_vett_1_14_port, g_vett_1_13_port, 
      g_vett_1_12_port, g_vett_1_11_port, g_vett_1_10_port, g_vett_1_9_port, 
      g_vett_1_8_port, g_vett_1_7_port, g_vett_1_6_port, g_vett_1_5_port, 
      g_vett_1_4_port, g_vett_1_3_port, g_vett_1_2_port, g_vett_1_1_port, 
      g_vett_1_0_port, g_vett_0_31_port, g_vett_0_30_port, g_vett_0_29_port, 
      g_vett_0_28_port, g_vett_0_27_port, g_vett_0_26_port, g_vett_0_25_port, 
      g_vett_0_24_port, g_vett_0_23_port, g_vett_0_22_port, g_vett_0_21_port, 
      g_vett_0_20_port, g_vett_0_19_port, g_vett_0_18_port, g_vett_0_17_port, 
      g_vett_0_16_port, g_vett_0_15_port, g_vett_0_14_port, g_vett_0_13_port, 
      g_vett_0_12_port, g_vett_0_11_port, g_vett_0_10_port, g_vett_0_9_port, 
      g_vett_0_8_port, g_vett_0_7_port, g_vett_0_6_port, g_vett_0_5_port, 
      g_vett_0_4_port, g_vett_0_3_port, g_vett_0_2_port, g_vett_0_1_port, 
      g_vett_0_0_port, n_1134 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Cin );
   
   PGblock_first : PG_block_0 port map( A => A(0), B => B(0), G => 
                           first_generate, P => p_vett_0_0_port);
   G_first : GENERAL_G_0 port map( G_in => first_generate, P_in => 
                           p_vett_0_0_port, G_in_prev => Cin, G_out => 
                           g_vett_0_0_port);
   PG_0_1 : PG_block_127 port map( A => A(1), B => B(1), G => g_vett_0_1_port, 
                           P => p_vett_0_1_port);
   PG_0_2 : PG_block_126 port map( A => A(2), B => B(2), G => g_vett_0_2_port, 
                           P => p_vett_0_2_port);
   PG_0_3 : PG_block_125 port map( A => A(3), B => B(3), G => g_vett_0_3_port, 
                           P => p_vett_0_3_port);
   PG_0_4 : PG_block_124 port map( A => A(4), B => B(4), G => g_vett_0_4_port, 
                           P => p_vett_0_4_port);
   PG_0_5 : PG_block_123 port map( A => A(5), B => B(5), G => g_vett_0_5_port, 
                           P => p_vett_0_5_port);
   PG_0_6 : PG_block_122 port map( A => A(6), B => B(6), G => g_vett_0_6_port, 
                           P => p_vett_0_6_port);
   PG_0_7 : PG_block_121 port map( A => A(7), B => B(7), G => g_vett_0_7_port, 
                           P => p_vett_0_7_port);
   PG_0_8 : PG_block_120 port map( A => A(8), B => B(8), G => g_vett_0_8_port, 
                           P => p_vett_0_8_port);
   PG_0_9 : PG_block_119 port map( A => A(9), B => B(9), G => g_vett_0_9_port, 
                           P => p_vett_0_9_port);
   PG_0_10 : PG_block_118 port map( A => A(10), B => B(10), G => 
                           g_vett_0_10_port, P => p_vett_0_10_port);
   PG_0_11 : PG_block_117 port map( A => A(11), B => B(11), G => 
                           g_vett_0_11_port, P => p_vett_0_11_port);
   PG_0_12 : PG_block_116 port map( A => A(12), B => B(12), G => 
                           g_vett_0_12_port, P => p_vett_0_12_port);
   PG_0_13 : PG_block_115 port map( A => A(13), B => B(13), G => 
                           g_vett_0_13_port, P => p_vett_0_13_port);
   PG_0_14 : PG_block_114 port map( A => A(14), B => B(14), G => 
                           g_vett_0_14_port, P => p_vett_0_14_port);
   PG_0_15 : PG_block_113 port map( A => A(15), B => B(15), G => 
                           g_vett_0_15_port, P => p_vett_0_15_port);
   PG_0_16 : PG_block_112 port map( A => A(16), B => B(16), G => 
                           g_vett_0_16_port, P => p_vett_0_16_port);
   PG_0_17 : PG_block_111 port map( A => A(17), B => B(17), G => 
                           g_vett_0_17_port, P => p_vett_0_17_port);
   PG_0_18 : PG_block_110 port map( A => A(18), B => B(18), G => 
                           g_vett_0_18_port, P => p_vett_0_18_port);
   PG_0_19 : PG_block_109 port map( A => A(19), B => B(19), G => 
                           g_vett_0_19_port, P => p_vett_0_19_port);
   PG_0_20 : PG_block_108 port map( A => A(20), B => B(20), G => 
                           g_vett_0_20_port, P => p_vett_0_20_port);
   PG_0_21 : PG_block_107 port map( A => A(21), B => B(21), G => 
                           g_vett_0_21_port, P => p_vett_0_21_port);
   PG_0_22 : PG_block_106 port map( A => A(22), B => B(22), G => 
                           g_vett_0_22_port, P => p_vett_0_22_port);
   PG_0_23 : PG_block_105 port map( A => A(23), B => B(23), G => 
                           g_vett_0_23_port, P => p_vett_0_23_port);
   PG_0_24 : PG_block_104 port map( A => A(24), B => B(24), G => 
                           g_vett_0_24_port, P => p_vett_0_24_port);
   PG_0_25 : PG_block_103 port map( A => A(25), B => B(25), G => 
                           g_vett_0_25_port, P => p_vett_0_25_port);
   PG_0_26 : PG_block_102 port map( A => A(26), B => B(26), G => 
                           g_vett_0_26_port, P => p_vett_0_26_port);
   PG_0_27 : PG_block_101 port map( A => A(27), B => B(27), G => 
                           g_vett_0_27_port, P => p_vett_0_27_port);
   PG_0_28 : PG_block_100 port map( A => A(28), B => B(28), G => 
                           g_vett_0_28_port, P => p_vett_0_28_port);
   PG_0_29 : PG_block_99 port map( A => A(29), B => B(29), G => 
                           g_vett_0_29_port, P => p_vett_0_29_port);
   PG_0_30 : PG_block_98 port map( A => A(30), B => B(30), G => 
                           g_vett_0_30_port, P => p_vett_0_30_port);
   PG_0_31 : PG_block_97 port map( A => A(31), B => B(31), G => 
                           g_vett_0_31_port, P => p_vett_0_31_port);
   G_0_0_0 : GENERAL_G_39 port map( G_in => g_vett_0_1_port, P_in => 
                           p_vett_0_1_port, G_in_prev => g_vett_0_0_port, G_out
                           => g_vett_1_0_port);
   PG_1_0_0 : GENERAL_PG_0 port map( G_in => g_vett_0_3_port, P_in => 
                           p_vett_0_3_port, G_in_prev => g_vett_0_2_port, 
                           P_in_prev => p_vett_0_2_port, G_out => 
                           g_vett_1_1_port, P_out => p_vett_1_1_port);
   G_1_0_0 : GENERAL_G_38 port map( G_in => g_vett_1_1_port, P_in => 
                           p_vett_1_1_port, G_in_prev => g_vett_1_0_port, G_out
                           => Co_1_port);
   PG_2_0_1 : GENERAL_PG_107 port map( G_in => g_vett_0_5_port, P_in => 
                           p_vett_0_5_port, G_in_prev => g_vett_0_4_port, 
                           P_in_prev => p_vett_0_4_port, G_out => 
                           g_vett_1_2_port, P_out => p_vett_1_2_port);
   PG_3_0_1 : GENERAL_PG_106 port map( G_in => g_vett_0_7_port, P_in => 
                           p_vett_0_7_port, G_in_prev => g_vett_0_6_port, 
                           P_in_prev => p_vett_0_6_port, G_out => 
                           g_vett_1_3_port, P_out => p_vett_1_3_port);
   PG_4_0_1 : GENERAL_PG_105 port map( G_in => g_vett_1_3_port, P_in => 
                           p_vett_1_3_port, G_in_prev => g_vett_1_2_port, 
                           P_in_prev => p_vett_1_2_port, G_out => 
                           g_vett_2_1_port, P_out => p_vett_2_1_port);
   PG_2_0_2 : GENERAL_PG_104 port map( G_in => g_vett_0_9_port, P_in => 
                           p_vett_0_9_port, G_in_prev => g_vett_0_8_port, 
                           P_in_prev => p_vett_0_8_port, G_out => 
                           g_vett_1_4_port, P_out => p_vett_1_4_port);
   PG_3_0_2 : GENERAL_PG_103 port map( G_in => g_vett_0_11_port, P_in => 
                           p_vett_0_11_port, G_in_prev => g_vett_0_10_port, 
                           P_in_prev => p_vett_0_10_port, G_out => 
                           g_vett_1_5_port, P_out => p_vett_1_5_port);
   PG_4_0_2 : GENERAL_PG_102 port map( G_in => g_vett_1_5_port, P_in => 
                           p_vett_1_5_port, G_in_prev => g_vett_1_4_port, 
                           P_in_prev => p_vett_1_4_port, G_out => 
                           g_vett_2_2_port, P_out => p_vett_2_2_port);
   PG_2_0_3 : GENERAL_PG_101 port map( G_in => g_vett_0_13_port, P_in => 
                           p_vett_0_13_port, G_in_prev => g_vett_0_12_port, 
                           P_in_prev => p_vett_0_12_port, G_out => 
                           g_vett_1_6_port, P_out => p_vett_1_6_port);
   PG_3_0_3 : GENERAL_PG_100 port map( G_in => g_vett_0_15_port, P_in => 
                           p_vett_0_15_port, G_in_prev => g_vett_0_14_port, 
                           P_in_prev => p_vett_0_14_port, G_out => 
                           g_vett_1_7_port, P_out => p_vett_1_7_port);
   PG_4_0_3 : GENERAL_PG_99 port map( G_in => g_vett_1_7_port, P_in => 
                           p_vett_1_7_port, G_in_prev => g_vett_1_6_port, 
                           P_in_prev => p_vett_1_6_port, G_out => 
                           g_vett_2_3_port, P_out => p_vett_2_3_port);
   PG_2_0_4 : GENERAL_PG_98 port map( G_in => g_vett_0_17_port, P_in => 
                           p_vett_0_17_port, G_in_prev => g_vett_0_16_port, 
                           P_in_prev => p_vett_0_16_port, G_out => 
                           g_vett_1_8_port, P_out => p_vett_1_8_port);
   PG_3_0_4 : GENERAL_PG_97 port map( G_in => g_vett_0_19_port, P_in => 
                           p_vett_0_19_port, G_in_prev => g_vett_0_18_port, 
                           P_in_prev => p_vett_0_18_port, G_out => 
                           g_vett_1_9_port, P_out => p_vett_1_9_port);
   PG_4_0_4 : GENERAL_PG_96 port map( G_in => g_vett_1_9_port, P_in => 
                           p_vett_1_9_port, G_in_prev => g_vett_1_8_port, 
                           P_in_prev => p_vett_1_8_port, G_out => 
                           g_vett_2_4_port, P_out => p_vett_2_4_port);
   PG_2_0_5 : GENERAL_PG_95 port map( G_in => g_vett_0_21_port, P_in => 
                           p_vett_0_21_port, G_in_prev => g_vett_0_20_port, 
                           P_in_prev => p_vett_0_20_port, G_out => 
                           g_vett_1_10_port, P_out => p_vett_1_10_port);
   PG_3_0_5 : GENERAL_PG_94 port map( G_in => g_vett_0_23_port, P_in => 
                           p_vett_0_23_port, G_in_prev => g_vett_0_22_port, 
                           P_in_prev => p_vett_0_22_port, G_out => 
                           g_vett_1_11_port, P_out => p_vett_1_11_port);
   PG_4_0_5 : GENERAL_PG_93 port map( G_in => g_vett_1_11_port, P_in => 
                           p_vett_1_11_port, G_in_prev => g_vett_1_10_port, 
                           P_in_prev => p_vett_1_10_port, G_out => 
                           g_vett_2_5_port, P_out => p_vett_2_5_port);
   PG_2_0_6 : GENERAL_PG_92 port map( G_in => g_vett_0_25_port, P_in => 
                           p_vett_0_25_port, G_in_prev => g_vett_0_24_port, 
                           P_in_prev => p_vett_0_24_port, G_out => 
                           g_vett_1_12_port, P_out => p_vett_1_12_port);
   PG_3_0_6 : GENERAL_PG_91 port map( G_in => g_vett_0_27_port, P_in => 
                           p_vett_0_27_port, G_in_prev => g_vett_0_26_port, 
                           P_in_prev => p_vett_0_26_port, G_out => 
                           g_vett_1_13_port, P_out => p_vett_1_13_port);
   PG_4_0_6 : GENERAL_PG_90 port map( G_in => g_vett_1_13_port, P_in => 
                           p_vett_1_13_port, G_in_prev => g_vett_1_12_port, 
                           P_in_prev => p_vett_1_12_port, G_out => 
                           g_vett_2_6_port, P_out => p_vett_2_6_port);
   PG_2_0_7 : GENERAL_PG_89 port map( G_in => g_vett_0_29_port, P_in => 
                           p_vett_0_29_port, G_in_prev => g_vett_0_28_port, 
                           P_in_prev => p_vett_0_28_port, G_out => 
                           g_vett_1_14_port, P_out => p_vett_1_14_port);
   PG_3_0_7 : GENERAL_PG_88 port map( G_in => g_vett_0_31_port, P_in => 
                           p_vett_0_31_port, G_in_prev => g_vett_0_30_port, 
                           P_in_prev => p_vett_0_30_port, G_out => 
                           g_vett_1_15_port, P_out => p_vett_1_15_port);
   PG_4_0_7 : GENERAL_PG_87 port map( G_in => g_vett_1_15_port, P_in => 
                           p_vett_1_15_port, G_in_prev => g_vett_1_14_port, 
                           P_in_prev => p_vett_1_14_port, G_out => 
                           g_vett_2_7_port, P_out => p_vett_2_7_port);
   G_2_1_0 : GENERAL_G_37 port map( G_in => g_vett_2_1_port, P_in => 
                           p_vett_2_1_port, G_in_prev => Co_1_port, G_out => 
                           Co_2_port);
   PG_5_1_0 : GENERAL_PG_86 port map( G_in => g_vett_2_3_port, P_in => 
                           p_vett_2_3_port, G_in_prev => g_vett_2_2_port, 
                           P_in_prev => p_vett_2_2_port, G_out => 
                           g_vett_3_1_port, P_out => p_vett_3_1_port);
   G_3_1_0 : GENERAL_G_36 port map( G_in => g_vett_2_2_port, P_in => 
                           p_vett_2_2_port, G_in_prev => Co_2_port, G_out => 
                           Co_3_port);
   G_4_1_0 : GENERAL_G_35 port map( G_in => g_vett_3_1_port, P_in => 
                           p_vett_3_1_port, G_in_prev => Co_2_port, G_out => 
                           Co_4_port);
   PG_6_1_1 : GENERAL_PG_85 port map( G_in => g_vett_2_5_port, P_in => 
                           p_vett_2_5_port, G_in_prev => g_vett_2_4_port, 
                           P_in_prev => p_vett_2_4_port, G_out => 
                           g_vett_3_2_port, P_out => p_vett_3_2_port);
   PG_7_1_1 : GENERAL_PG_84 port map( G_in => g_vett_2_7_port, P_in => 
                           p_vett_2_7_port, G_in_prev => g_vett_2_6_port, 
                           P_in_prev => p_vett_2_6_port, G_out => 
                           g_vett_3_3_port, P_out => p_vett_3_3_port);
   PG_8_1_1 : GENERAL_PG_83 port map( G_in => g_vett_2_6_port, P_in => 
                           p_vett_2_6_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_2_port, P_out => p_vett_4_2_port);
   PG_9_1_1 : GENERAL_PG_82 port map( G_in => g_vett_3_3_port, P_in => 
                           p_vett_3_3_port, G_in_prev => g_vett_3_2_port, 
                           P_in_prev => p_vett_3_2_port, G_out => 
                           g_vett_4_3_port, P_out => p_vett_4_3_port);
   G_5_2_0 : GENERAL_G_34 port map( G_in => g_vett_2_4_port, P_in => 
                           p_vett_2_4_port, G_in_prev => Co_4_port, G_out => 
                           Co_5_port);
   G_6_2_1 : GENERAL_G_33 port map( G_in => g_vett_3_2_port, P_in => 
                           p_vett_3_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_6_port);
   G_7_2_2 : GENERAL_G_32 port map( G_in => g_vett_4_2_port, P_in => 
                           p_vett_4_2_port, G_in_prev => Co_4_port, G_out => 
                           Co_7_port);
   G_8_2_3 : GENERAL_G_31 port map( G_in => g_vett_4_3_port, P_in => 
                           p_vett_4_3_port, G_in_prev => Co_4_port, G_out => 
                           n_1134);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n78, ZN => n68);
   U2 : INV_X1 port map( A => n78, ZN => n69);
   U3 : BUF_X1 port map( A => n33, Z => n70);
   U4 : BUF_X1 port map( A => n67, Z => n76);
   U5 : BUF_X1 port map( A => n66, Z => n75);
   U6 : BUF_X1 port map( A => n66, Z => n73);
   U7 : BUF_X1 port map( A => n33, Z => n72);
   U8 : BUF_X1 port map( A => n66, Z => n74);
   U9 : BUF_X1 port map( A => n33, Z => n71);
   U10 : BUF_X1 port map( A => n67, Z => n78);
   U11 : BUF_X1 port map( A => n67, Z => n77);
   U12 : BUF_X1 port map( A => SEL, Z => n67);
   U13 : BUF_X1 port map( A => SEL, Z => n66);
   U14 : BUF_X1 port map( A => SEL, Z => n33);
   U15 : INV_X1 port map( A => n136, ZN => Y(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n68, B1 => B(3), B2 => n71, ZN =>
                           n136);
   U17 : INV_X1 port map( A => n137, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n69, B1 => B(4), B2 => n71, ZN =>
                           n137);
   U19 : INV_X1 port map( A => n138, ZN => Y(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n68, B1 => B(5), B2 => n70, ZN =>
                           n138);
   U21 : INV_X1 port map( A => n139, ZN => Y(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n69, B1 => B(6), B2 => n70, ZN =>
                           n139);
   U23 : INV_X1 port map( A => n140, ZN => Y(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n68, B1 => B(7), B2 => n70, ZN =>
                           n140);
   U25 : INV_X1 port map( A => n141, ZN => Y(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n69, B1 => B(8), B2 => n70, ZN =>
                           n141);
   U27 : INV_X1 port map( A => n142, ZN => Y(9));
   U28 : AOI22_X1 port map( A1 => A(9), A2 => n68, B1 => n77, B2 => B(9), ZN =>
                           n142);
   U29 : INV_X1 port map( A => n135, ZN => Y(31));
   U30 : AOI22_X1 port map( A1 => A(31), A2 => n69, B1 => B(31), B2 => n71, ZN 
                           => n135);
   U31 : INV_X1 port map( A => n111, ZN => Y(0));
   U32 : AOI22_X1 port map( A1 => A(0), A2 => n68, B1 => B(0), B2 => n77, ZN =>
                           n111);
   U33 : INV_X1 port map( A => n122, ZN => Y(1));
   U34 : AOI22_X1 port map( A1 => A(1), A2 => n68, B1 => B(1), B2 => n74, ZN =>
                           n122);
   U35 : INV_X1 port map( A => n133, ZN => Y(2));
   U36 : AOI22_X1 port map( A1 => A(2), A2 => n69, B1 => B(2), B2 => n71, ZN =>
                           n133);
   U37 : INV_X1 port map( A => n112, ZN => Y(10));
   U38 : AOI22_X1 port map( A1 => A(10), A2 => n68, B1 => B(10), B2 => n77, ZN 
                           => n112);
   U39 : INV_X1 port map( A => n113, ZN => Y(11));
   U40 : AOI22_X1 port map( A1 => A(11), A2 => n68, B1 => B(11), B2 => n77, ZN 
                           => n113);
   U41 : INV_X1 port map( A => n114, ZN => Y(12));
   U42 : AOI22_X1 port map( A1 => A(12), A2 => n68, B1 => B(12), B2 => n76, ZN 
                           => n114);
   U43 : INV_X1 port map( A => n115, ZN => Y(13));
   U44 : AOI22_X1 port map( A1 => A(13), A2 => n68, B1 => B(13), B2 => n76, ZN 
                           => n115);
   U45 : INV_X1 port map( A => n116, ZN => Y(14));
   U46 : AOI22_X1 port map( A1 => A(14), A2 => n68, B1 => B(14), B2 => n76, ZN 
                           => n116);
   U47 : INV_X1 port map( A => n117, ZN => Y(15));
   U48 : AOI22_X1 port map( A1 => A(15), A2 => n68, B1 => B(15), B2 => n76, ZN 
                           => n117);
   U49 : INV_X1 port map( A => n118, ZN => Y(16));
   U50 : AOI22_X1 port map( A1 => A(16), A2 => n68, B1 => B(16), B2 => n75, ZN 
                           => n118);
   U51 : INV_X1 port map( A => n119, ZN => Y(17));
   U52 : AOI22_X1 port map( A1 => A(17), A2 => n68, B1 => B(17), B2 => n75, ZN 
                           => n119);
   U53 : INV_X1 port map( A => n120, ZN => Y(18));
   U54 : AOI22_X1 port map( A1 => A(18), A2 => n68, B1 => B(18), B2 => n75, ZN 
                           => n120);
   U55 : INV_X1 port map( A => n121, ZN => Y(19));
   U56 : AOI22_X1 port map( A1 => A(19), A2 => n68, B1 => B(19), B2 => n75, ZN 
                           => n121);
   U57 : INV_X1 port map( A => n123, ZN => Y(20));
   U58 : AOI22_X1 port map( A1 => A(20), A2 => n69, B1 => B(20), B2 => n74, ZN 
                           => n123);
   U59 : INV_X1 port map( A => n124, ZN => Y(21));
   U60 : AOI22_X1 port map( A1 => A(21), A2 => n69, B1 => B(21), B2 => n74, ZN 
                           => n124);
   U61 : INV_X1 port map( A => n125, ZN => Y(22));
   U62 : AOI22_X1 port map( A1 => A(22), A2 => n69, B1 => B(22), B2 => n73, ZN 
                           => n125);
   U63 : INV_X1 port map( A => n126, ZN => Y(23));
   U64 : AOI22_X1 port map( A1 => A(23), A2 => n69, B1 => B(23), B2 => n73, ZN 
                           => n126);
   U65 : INV_X1 port map( A => n127, ZN => Y(24));
   U66 : AOI22_X1 port map( A1 => A(24), A2 => n69, B1 => B(24), B2 => n73, ZN 
                           => n127);
   U67 : INV_X1 port map( A => n128, ZN => Y(25));
   U68 : AOI22_X1 port map( A1 => A(25), A2 => n69, B1 => B(25), B2 => n73, ZN 
                           => n128);
   U69 : INV_X1 port map( A => n129, ZN => Y(26));
   U70 : AOI22_X1 port map( A1 => A(26), A2 => n69, B1 => B(26), B2 => n72, ZN 
                           => n129);
   U71 : INV_X1 port map( A => n130, ZN => Y(27));
   U72 : AOI22_X1 port map( A1 => A(27), A2 => n69, B1 => B(27), B2 => n72, ZN 
                           => n130);
   U73 : INV_X1 port map( A => n131, ZN => Y(28));
   U74 : AOI22_X1 port map( A1 => A(28), A2 => n69, B1 => B(28), B2 => n72, ZN 
                           => n131);
   U75 : INV_X1 port map( A => n132, ZN => Y(29));
   U76 : AOI22_X1 port map( A1 => A(29), A2 => n69, B1 => B(29), B2 => n72, ZN 
                           => n132);
   U77 : INV_X1 port map( A => n134, ZN => Y(30));
   U78 : AOI22_X1 port map( A1 => A(30), A2 => n69, B1 => B(30), B2 => n74, ZN 
                           => n134);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_1 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_1;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42
      , n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n47, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n49, Q => Q(30), 
                           QN => n67);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n49, Q => Q(29), 
                           QN => n68);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n49, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n49, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n48, Q => Q(26), 
                           QN => n71);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n49, Q => Q(25), 
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n48, Q => Q(24), 
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n48, Q => Q(23), 
                           QN => n74);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n48, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n48, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n49, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n48, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n48, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n49, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n48, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n48, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n48, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n47, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n48, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n47, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n47, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n47, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n47, Q => Q(8), 
                           QN => n89);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n47, Q => Q(7), 
                           QN => n90);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n47, Q => Q(6), 
                           QN => n91);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n47, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n47, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n47, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n47, Q => Q(2), 
                           QN => n95);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n48, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n49, Q => Q(0), 
                           QN => n97);
   U2 : INV_X1 port map( A => n46, ZN => n37);
   U3 : INV_X1 port map( A => n46, ZN => n36);
   U4 : BUF_X1 port map( A => n35, Z => n46);
   U5 : BUF_X1 port map( A => n34, Z => n41);
   U6 : BUF_X1 port map( A => n34, Z => n42);
   U7 : BUF_X1 port map( A => n35, Z => n44);
   U8 : BUF_X1 port map( A => n33, Z => n38);
   U9 : BUF_X1 port map( A => n33, Z => n39);
   U10 : BUF_X1 port map( A => n33, Z => n40);
   U11 : BUF_X1 port map( A => n34, Z => n43);
   U12 : BUF_X1 port map( A => n35, Z => n45);
   U13 : BUF_X1 port map( A => RESET_n, Z => n48);
   U14 : BUF_X1 port map( A => RESET_n, Z => n47);
   U15 : BUF_X1 port map( A => RESET_n, Z => n49);
   U16 : BUF_X1 port map( A => Enable_n, Z => n35);
   U17 : BUF_X1 port map( A => Enable_n, Z => n33);
   U18 : BUF_X1 port map( A => Enable_n, Z => n34);
   U19 : OAI22_X1 port map( A1 => n70, A2 => n37, B1 => n39, B2 => n54, ZN => 
                           n5);
   U20 : INV_X1 port map( A => D(27), ZN => n54);
   U21 : OAI22_X1 port map( A1 => n69, A2 => n36, B1 => n39, B2 => n53, ZN => 
                           n4);
   U22 : INV_X1 port map( A => D(28), ZN => n53);
   U23 : OAI22_X1 port map( A1 => n97, A2 => n37, B1 => n39, B2 => n113, ZN => 
                           n32);
   U24 : INV_X1 port map( A => D(0), ZN => n113);
   U25 : OAI22_X1 port map( A1 => n96, A2 => n36, B1 => n39, B2 => n112, ZN => 
                           n31);
   U26 : INV_X1 port map( A => D(1), ZN => n112);
   U27 : OAI22_X1 port map( A1 => n74, A2 => n37, B1 => n38, B2 => n58, ZN => 
                           n9);
   U28 : INV_X1 port map( A => D(23), ZN => n58);
   U29 : OAI22_X1 port map( A1 => n73, A2 => n36, B1 => n38, B2 => n57, ZN => 
                           n8);
   U30 : INV_X1 port map( A => D(24), ZN => n57);
   U31 : OAI22_X1 port map( A1 => n72, A2 => n37, B1 => n38, B2 => n56, ZN => 
                           n7);
   U32 : INV_X1 port map( A => D(25), ZN => n56);
   U33 : OAI22_X1 port map( A1 => n71, A2 => n36, B1 => n38, B2 => n55, ZN => 
                           n6);
   U34 : INV_X1 port map( A => D(26), ZN => n55);
   U35 : OAI22_X1 port map( A1 => n95, A2 => n37, B1 => n40, B2 => n111, ZN => 
                           n30);
   U36 : INV_X1 port map( A => D(2), ZN => n111);
   U37 : OAI22_X1 port map( A1 => n94, A2 => n37, B1 => n40, B2 => n110, ZN => 
                           n29);
   U38 : INV_X1 port map( A => D(3), ZN => n110);
   U39 : OAI22_X1 port map( A1 => n93, A2 => n37, B1 => n40, B2 => n109, ZN => 
                           n28);
   U40 : INV_X1 port map( A => D(4), ZN => n109);
   U41 : OAI22_X1 port map( A1 => n92, A2 => n37, B1 => n41, B2 => n108, ZN => 
                           n27);
   U42 : INV_X1 port map( A => D(5), ZN => n108);
   U43 : OAI22_X1 port map( A1 => n91, A2 => n37, B1 => n41, B2 => n107, ZN => 
                           n26);
   U44 : INV_X1 port map( A => D(6), ZN => n107);
   U45 : OAI22_X1 port map( A1 => n90, A2 => n37, B1 => n41, B2 => n106, ZN => 
                           n25);
   U46 : INV_X1 port map( A => D(7), ZN => n106);
   U47 : OAI22_X1 port map( A1 => n89, A2 => n37, B1 => n41, B2 => n105, ZN => 
                           n24);
   U48 : INV_X1 port map( A => D(8), ZN => n105);
   U49 : OAI22_X1 port map( A1 => n88, A2 => n37, B1 => n42, B2 => n104, ZN => 
                           n23);
   U50 : INV_X1 port map( A => D(9), ZN => n104);
   U51 : OAI22_X1 port map( A1 => n87, A2 => n37, B1 => n42, B2 => n103, ZN => 
                           n22);
   U52 : INV_X1 port map( A => D(10), ZN => n103);
   U53 : OAI22_X1 port map( A1 => n86, A2 => n37, B1 => n42, B2 => n102, ZN => 
                           n21);
   U54 : INV_X1 port map( A => D(11), ZN => n102);
   U55 : OAI22_X1 port map( A1 => n85, A2 => n37, B1 => n42, B2 => n101, ZN => 
                           n20);
   U56 : INV_X1 port map( A => D(12), ZN => n101);
   U57 : OAI22_X1 port map( A1 => n84, A2 => n36, B1 => n43, B2 => n100, ZN => 
                           n19);
   U58 : INV_X1 port map( A => D(13), ZN => n100);
   U59 : OAI22_X1 port map( A1 => n83, A2 => n36, B1 => n43, B2 => n99, ZN => 
                           n18);
   U60 : INV_X1 port map( A => D(14), ZN => n99);
   U61 : OAI22_X1 port map( A1 => n82, A2 => n36, B1 => n43, B2 => n98, ZN => 
                           n17);
   U62 : INV_X1 port map( A => D(15), ZN => n98);
   U63 : OAI22_X1 port map( A1 => n81, A2 => n36, B1 => n44, B2 => n65, ZN => 
                           n16);
   U64 : INV_X1 port map( A => D(16), ZN => n65);
   U65 : OAI22_X1 port map( A1 => n80, A2 => n36, B1 => n44, B2 => n64, ZN => 
                           n15);
   U66 : INV_X1 port map( A => D(17), ZN => n64);
   U67 : OAI22_X1 port map( A1 => n79, A2 => n36, B1 => n44, B2 => n63, ZN => 
                           n14);
   U68 : INV_X1 port map( A => D(18), ZN => n63);
   U69 : OAI22_X1 port map( A1 => n78, A2 => n36, B1 => n44, B2 => n62, ZN => 
                           n13);
   U70 : INV_X1 port map( A => D(19), ZN => n62);
   U71 : OAI22_X1 port map( A1 => n77, A2 => n36, B1 => n45, B2 => n61, ZN => 
                           n12);
   U72 : INV_X1 port map( A => D(20), ZN => n61);
   U73 : OAI22_X1 port map( A1 => n76, A2 => n36, B1 => n45, B2 => n60, ZN => 
                           n11);
   U74 : INV_X1 port map( A => D(21), ZN => n60);
   U75 : OAI22_X1 port map( A1 => n75, A2 => n36, B1 => n45, B2 => n59, ZN => 
                           n10);
   U76 : INV_X1 port map( A => D(22), ZN => n59);
   U77 : OAI22_X1 port map( A1 => n68, A2 => n37, B1 => n40, B2 => n52, ZN => 
                           n3);
   U78 : INV_X1 port map( A => D(29), ZN => n52);
   U79 : OAI22_X1 port map( A1 => n67, A2 => n36, B1 => n43, B2 => n51, ZN => 
                           n2);
   U80 : INV_X1 port map( A => D(30), ZN => n51);
   U81 : OAI22_X1 port map( A1 => n66, A2 => n36, B1 => n45, B2 => n50, ZN => 
                           n1);
   U82 : INV_X1 port map( A => D(31), ZN => n50);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_2 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_2;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n49, Q => Q(31), 
                           QN => n145);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n49, Q => Q(30), 
                           QN => n144);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n49, Q => Q(29), 
                           QN => n143);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n49, Q => Q(28), 
                           QN => n142);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n49, Q => Q(27), 
                           QN => n141);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n49, Q => Q(26), 
                           QN => n140);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n49, Q => Q(25), 
                           QN => n139);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n49, Q => Q(24), 
                           QN => n138);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n48, Q => Q(23), 
                           QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n48, Q => Q(22),
                           QN => n136);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n48, Q => Q(21),
                           QN => n135);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n48, Q => Q(20),
                           QN => n134);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n48, Q => Q(19),
                           QN => n133);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n48, Q => Q(18),
                           QN => n132);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n48, Q => Q(17),
                           QN => n131);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n48, Q => Q(16),
                           QN => n130);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n48, Q => Q(15),
                           QN => n129);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n48, Q => Q(14),
                           QN => n128);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n48, Q => Q(13),
                           QN => n127);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n48, Q => Q(12),
                           QN => n126);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n47, Q => Q(11),
                           QN => n125);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n47, Q => Q(10),
                           QN => n124);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n47, Q => Q(9), 
                           QN => n123);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n47, Q => Q(8), 
                           QN => n122);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n47, Q => Q(7), 
                           QN => n121);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n47, Q => Q(6), 
                           QN => n120);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n47, Q => Q(5), 
                           QN => n119);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n47, Q => Q(4), 
                           QN => n118);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n47, Q => Q(3), 
                           QN => n117);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n47, Q => Q(2), 
                           QN => n116);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n47, Q => Q(1), 
                           QN => n115);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n47, Q => Q(0), 
                           QN => n114);
   U2 : INV_X1 port map( A => n46, ZN => n37);
   U3 : INV_X1 port map( A => n46, ZN => n36);
   U4 : BUF_X1 port map( A => n35, Z => n46);
   U5 : BUF_X1 port map( A => n34, Z => n41);
   U6 : BUF_X1 port map( A => n34, Z => n42);
   U7 : BUF_X1 port map( A => n35, Z => n44);
   U8 : BUF_X1 port map( A => n33, Z => n38);
   U9 : BUF_X1 port map( A => n33, Z => n39);
   U10 : BUF_X1 port map( A => n33, Z => n40);
   U11 : BUF_X1 port map( A => n34, Z => n43);
   U12 : BUF_X1 port map( A => n35, Z => n45);
   U13 : BUF_X1 port map( A => RESET_n, Z => n47);
   U14 : BUF_X1 port map( A => RESET_n, Z => n48);
   U15 : BUF_X1 port map( A => RESET_n, Z => n49);
   U16 : BUF_X1 port map( A => Enable_n, Z => n35);
   U17 : BUF_X1 port map( A => Enable_n, Z => n33);
   U18 : BUF_X1 port map( A => Enable_n, Z => n34);
   U19 : OAI22_X1 port map( A1 => n114, A2 => n37, B1 => n39, B2 => n113, ZN =>
                           n32);
   U20 : INV_X1 port map( A => D(0), ZN => n113);
   U21 : OAI22_X1 port map( A1 => n115, A2 => n36, B1 => n39, B2 => n112, ZN =>
                           n31);
   U22 : INV_X1 port map( A => D(1), ZN => n112);
   U23 : OAI22_X1 port map( A1 => n137, A2 => n37, B1 => n38, B2 => n58, ZN => 
                           n9);
   U24 : INV_X1 port map( A => D(23), ZN => n58);
   U25 : OAI22_X1 port map( A1 => n138, A2 => n36, B1 => n38, B2 => n57, ZN => 
                           n8);
   U26 : INV_X1 port map( A => D(24), ZN => n57);
   U27 : OAI22_X1 port map( A1 => n139, A2 => n37, B1 => n38, B2 => n56, ZN => 
                           n7);
   U28 : INV_X1 port map( A => D(25), ZN => n56);
   U29 : OAI22_X1 port map( A1 => n140, A2 => n36, B1 => n38, B2 => n55, ZN => 
                           n6);
   U30 : INV_X1 port map( A => D(26), ZN => n55);
   U31 : OAI22_X1 port map( A1 => n141, A2 => n37, B1 => n39, B2 => n54, ZN => 
                           n5);
   U32 : INV_X1 port map( A => D(27), ZN => n54);
   U33 : OAI22_X1 port map( A1 => n142, A2 => n36, B1 => n39, B2 => n53, ZN => 
                           n4);
   U34 : INV_X1 port map( A => D(28), ZN => n53);
   U35 : OAI22_X1 port map( A1 => n116, A2 => n37, B1 => n40, B2 => n111, ZN =>
                           n30);
   U36 : INV_X1 port map( A => D(2), ZN => n111);
   U37 : OAI22_X1 port map( A1 => n117, A2 => n37, B1 => n40, B2 => n110, ZN =>
                           n29);
   U38 : INV_X1 port map( A => D(3), ZN => n110);
   U39 : OAI22_X1 port map( A1 => n118, A2 => n37, B1 => n40, B2 => n109, ZN =>
                           n28);
   U40 : INV_X1 port map( A => D(4), ZN => n109);
   U41 : OAI22_X1 port map( A1 => n119, A2 => n37, B1 => n41, B2 => n108, ZN =>
                           n27);
   U42 : INV_X1 port map( A => D(5), ZN => n108);
   U43 : OAI22_X1 port map( A1 => n120, A2 => n37, B1 => n41, B2 => n107, ZN =>
                           n26);
   U44 : INV_X1 port map( A => D(6), ZN => n107);
   U45 : OAI22_X1 port map( A1 => n121, A2 => n37, B1 => n41, B2 => n106, ZN =>
                           n25);
   U46 : INV_X1 port map( A => D(7), ZN => n106);
   U47 : OAI22_X1 port map( A1 => n122, A2 => n37, B1 => n41, B2 => n105, ZN =>
                           n24);
   U48 : INV_X1 port map( A => D(8), ZN => n105);
   U49 : OAI22_X1 port map( A1 => n123, A2 => n37, B1 => n42, B2 => n104, ZN =>
                           n23);
   U50 : INV_X1 port map( A => D(9), ZN => n104);
   U51 : OAI22_X1 port map( A1 => n124, A2 => n37, B1 => n42, B2 => n103, ZN =>
                           n22);
   U52 : INV_X1 port map( A => D(10), ZN => n103);
   U53 : OAI22_X1 port map( A1 => n125, A2 => n37, B1 => n42, B2 => n102, ZN =>
                           n21);
   U54 : INV_X1 port map( A => D(11), ZN => n102);
   U55 : OAI22_X1 port map( A1 => n126, A2 => n37, B1 => n42, B2 => n101, ZN =>
                           n20);
   U56 : INV_X1 port map( A => D(12), ZN => n101);
   U57 : OAI22_X1 port map( A1 => n127, A2 => n36, B1 => n43, B2 => n100, ZN =>
                           n19);
   U58 : INV_X1 port map( A => D(13), ZN => n100);
   U59 : OAI22_X1 port map( A1 => n128, A2 => n36, B1 => n43, B2 => n99, ZN => 
                           n18);
   U60 : INV_X1 port map( A => D(14), ZN => n99);
   U61 : OAI22_X1 port map( A1 => n129, A2 => n36, B1 => n43, B2 => n98, ZN => 
                           n17);
   U62 : INV_X1 port map( A => D(15), ZN => n98);
   U63 : OAI22_X1 port map( A1 => n130, A2 => n36, B1 => n44, B2 => n65, ZN => 
                           n16);
   U64 : INV_X1 port map( A => D(16), ZN => n65);
   U65 : OAI22_X1 port map( A1 => n131, A2 => n36, B1 => n44, B2 => n64, ZN => 
                           n15);
   U66 : INV_X1 port map( A => D(17), ZN => n64);
   U67 : OAI22_X1 port map( A1 => n132, A2 => n36, B1 => n44, B2 => n63, ZN => 
                           n14);
   U68 : INV_X1 port map( A => D(18), ZN => n63);
   U69 : OAI22_X1 port map( A1 => n133, A2 => n36, B1 => n44, B2 => n62, ZN => 
                           n13);
   U70 : INV_X1 port map( A => D(19), ZN => n62);
   U71 : OAI22_X1 port map( A1 => n134, A2 => n36, B1 => n45, B2 => n61, ZN => 
                           n12);
   U72 : INV_X1 port map( A => D(20), ZN => n61);
   U73 : OAI22_X1 port map( A1 => n135, A2 => n36, B1 => n45, B2 => n60, ZN => 
                           n11);
   U74 : INV_X1 port map( A => D(21), ZN => n60);
   U75 : OAI22_X1 port map( A1 => n136, A2 => n36, B1 => n45, B2 => n59, ZN => 
                           n10);
   U76 : INV_X1 port map( A => D(22), ZN => n59);
   U77 : OAI22_X1 port map( A1 => n143, A2 => n37, B1 => n40, B2 => n52, ZN => 
                           n3);
   U78 : INV_X1 port map( A => D(29), ZN => n52);
   U79 : OAI22_X1 port map( A1 => n144, A2 => n36, B1 => n43, B2 => n51, ZN => 
                           n2);
   U80 : INV_X1 port map( A => D(30), ZN => n51);
   U81 : OAI22_X1 port map( A1 => n145, A2 => n36, B1 => n45, B2 => n50, ZN => 
                           n1);
   U82 : INV_X1 port map( A => D(31), ZN => n50);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_3 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_3;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n47, Q => Q(31), 
                           QN => n145);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n47, Q => Q(30), 
                           QN => n144);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n47, Q => Q(29), 
                           QN => n143);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n47, Q => Q(28), 
                           QN => n142);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n47, Q => Q(27), 
                           QN => n141);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n47, Q => Q(26), 
                           QN => n140);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n47, Q => Q(25), 
                           QN => n139);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n47, Q => Q(24), 
                           QN => n138);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n47, Q => Q(23), 
                           QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n47, Q => Q(22),
                           QN => n136);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n47, Q => Q(21),
                           QN => n135);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n47, Q => Q(20),
                           QN => n134);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n48, Q => Q(19),
                           QN => n133);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n48, Q => Q(18),
                           QN => n132);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n48, Q => Q(17),
                           QN => n131);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n48, Q => Q(16),
                           QN => n130);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n48, Q => Q(15),
                           QN => n129);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n48, Q => Q(14),
                           QN => n128);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n48, Q => Q(13),
                           QN => n127);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n48, Q => Q(12),
                           QN => n126);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n48, Q => Q(11),
                           QN => n125);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n48, Q => Q(10),
                           QN => n124);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n48, Q => Q(9), 
                           QN => n123);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n48, Q => Q(8), 
                           QN => n122);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n49, Q => Q(7), 
                           QN => n121);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n49, Q => Q(6), 
                           QN => n120);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n49, Q => Q(5), 
                           QN => n119);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n49, Q => Q(4), 
                           QN => n118);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n49, Q => Q(3), 
                           QN => n117);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n49, Q => Q(2), 
                           QN => n116);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n49, Q => Q(1), 
                           QN => n115);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n49, Q => Q(0), 
                           QN => n114);
   U2 : INV_X1 port map( A => n46, ZN => n37);
   U3 : INV_X1 port map( A => n46, ZN => n36);
   U4 : BUF_X1 port map( A => n35, Z => n46);
   U5 : BUF_X1 port map( A => n34, Z => n41);
   U6 : BUF_X1 port map( A => n34, Z => n42);
   U7 : BUF_X1 port map( A => n35, Z => n44);
   U8 : BUF_X1 port map( A => n33, Z => n38);
   U9 : BUF_X1 port map( A => n33, Z => n39);
   U10 : BUF_X1 port map( A => n33, Z => n40);
   U11 : BUF_X1 port map( A => n34, Z => n43);
   U12 : BUF_X1 port map( A => n35, Z => n45);
   U13 : BUF_X1 port map( A => RESET_n, Z => n48);
   U14 : BUF_X1 port map( A => RESET_n, Z => n47);
   U15 : BUF_X1 port map( A => RESET_n, Z => n49);
   U16 : BUF_X1 port map( A => Enable_n, Z => n35);
   U17 : BUF_X1 port map( A => Enable_n, Z => n33);
   U18 : BUF_X1 port map( A => Enable_n, Z => n34);
   U19 : OAI22_X1 port map( A1 => n114, A2 => n37, B1 => n39, B2 => n113, ZN =>
                           n32);
   U20 : INV_X1 port map( A => D(0), ZN => n113);
   U21 : OAI22_X1 port map( A1 => n115, A2 => n36, B1 => n39, B2 => n112, ZN =>
                           n31);
   U22 : INV_X1 port map( A => D(1), ZN => n112);
   U23 : OAI22_X1 port map( A1 => n137, A2 => n37, B1 => n38, B2 => n58, ZN => 
                           n9);
   U24 : INV_X1 port map( A => D(23), ZN => n58);
   U25 : OAI22_X1 port map( A1 => n138, A2 => n36, B1 => n38, B2 => n57, ZN => 
                           n8);
   U26 : INV_X1 port map( A => D(24), ZN => n57);
   U27 : OAI22_X1 port map( A1 => n139, A2 => n37, B1 => n38, B2 => n56, ZN => 
                           n7);
   U28 : INV_X1 port map( A => D(25), ZN => n56);
   U29 : OAI22_X1 port map( A1 => n140, A2 => n36, B1 => n38, B2 => n55, ZN => 
                           n6);
   U30 : INV_X1 port map( A => D(26), ZN => n55);
   U31 : OAI22_X1 port map( A1 => n141, A2 => n37, B1 => n39, B2 => n54, ZN => 
                           n5);
   U32 : INV_X1 port map( A => D(27), ZN => n54);
   U33 : OAI22_X1 port map( A1 => n142, A2 => n36, B1 => n39, B2 => n53, ZN => 
                           n4);
   U34 : INV_X1 port map( A => D(28), ZN => n53);
   U35 : OAI22_X1 port map( A1 => n116, A2 => n37, B1 => n40, B2 => n111, ZN =>
                           n30);
   U36 : INV_X1 port map( A => D(2), ZN => n111);
   U37 : OAI22_X1 port map( A1 => n117, A2 => n37, B1 => n40, B2 => n110, ZN =>
                           n29);
   U38 : INV_X1 port map( A => D(3), ZN => n110);
   U39 : OAI22_X1 port map( A1 => n118, A2 => n37, B1 => n40, B2 => n109, ZN =>
                           n28);
   U40 : INV_X1 port map( A => D(4), ZN => n109);
   U41 : OAI22_X1 port map( A1 => n119, A2 => n37, B1 => n41, B2 => n108, ZN =>
                           n27);
   U42 : INV_X1 port map( A => D(5), ZN => n108);
   U43 : OAI22_X1 port map( A1 => n120, A2 => n37, B1 => n41, B2 => n107, ZN =>
                           n26);
   U44 : INV_X1 port map( A => D(6), ZN => n107);
   U45 : OAI22_X1 port map( A1 => n121, A2 => n37, B1 => n41, B2 => n106, ZN =>
                           n25);
   U46 : INV_X1 port map( A => D(7), ZN => n106);
   U47 : OAI22_X1 port map( A1 => n122, A2 => n37, B1 => n41, B2 => n105, ZN =>
                           n24);
   U48 : INV_X1 port map( A => D(8), ZN => n105);
   U49 : OAI22_X1 port map( A1 => n123, A2 => n37, B1 => n42, B2 => n104, ZN =>
                           n23);
   U50 : INV_X1 port map( A => D(9), ZN => n104);
   U51 : OAI22_X1 port map( A1 => n124, A2 => n37, B1 => n42, B2 => n103, ZN =>
                           n22);
   U52 : INV_X1 port map( A => D(10), ZN => n103);
   U53 : OAI22_X1 port map( A1 => n125, A2 => n37, B1 => n42, B2 => n102, ZN =>
                           n21);
   U54 : INV_X1 port map( A => D(11), ZN => n102);
   U55 : OAI22_X1 port map( A1 => n126, A2 => n37, B1 => n42, B2 => n101, ZN =>
                           n20);
   U56 : INV_X1 port map( A => D(12), ZN => n101);
   U57 : OAI22_X1 port map( A1 => n127, A2 => n36, B1 => n43, B2 => n100, ZN =>
                           n19);
   U58 : INV_X1 port map( A => D(13), ZN => n100);
   U59 : OAI22_X1 port map( A1 => n128, A2 => n36, B1 => n43, B2 => n99, ZN => 
                           n18);
   U60 : INV_X1 port map( A => D(14), ZN => n99);
   U61 : OAI22_X1 port map( A1 => n129, A2 => n36, B1 => n43, B2 => n98, ZN => 
                           n17);
   U62 : INV_X1 port map( A => D(15), ZN => n98);
   U63 : OAI22_X1 port map( A1 => n130, A2 => n36, B1 => n44, B2 => n65, ZN => 
                           n16);
   U64 : INV_X1 port map( A => D(16), ZN => n65);
   U65 : OAI22_X1 port map( A1 => n131, A2 => n36, B1 => n44, B2 => n64, ZN => 
                           n15);
   U66 : INV_X1 port map( A => D(17), ZN => n64);
   U67 : OAI22_X1 port map( A1 => n132, A2 => n36, B1 => n44, B2 => n63, ZN => 
                           n14);
   U68 : INV_X1 port map( A => D(18), ZN => n63);
   U69 : OAI22_X1 port map( A1 => n133, A2 => n36, B1 => n44, B2 => n62, ZN => 
                           n13);
   U70 : INV_X1 port map( A => D(19), ZN => n62);
   U71 : OAI22_X1 port map( A1 => n134, A2 => n36, B1 => n45, B2 => n61, ZN => 
                           n12);
   U72 : INV_X1 port map( A => D(20), ZN => n61);
   U73 : OAI22_X1 port map( A1 => n135, A2 => n36, B1 => n45, B2 => n60, ZN => 
                           n11);
   U74 : INV_X1 port map( A => D(21), ZN => n60);
   U75 : OAI22_X1 port map( A1 => n136, A2 => n36, B1 => n45, B2 => n59, ZN => 
                           n10);
   U76 : INV_X1 port map( A => D(22), ZN => n59);
   U77 : OAI22_X1 port map( A1 => n143, A2 => n37, B1 => n40, B2 => n52, ZN => 
                           n3);
   U78 : INV_X1 port map( A => D(29), ZN => n52);
   U79 : OAI22_X1 port map( A1 => n144, A2 => n36, B1 => n43, B2 => n51, ZN => 
                           n2);
   U80 : INV_X1 port map( A => D(30), ZN => n51);
   U81 : OAI22_X1 port map( A1 => n145, A2 => n36, B1 => n45, B2 => n50, ZN => 
                           n1);
   U82 : INV_X1 port map( A => D(31), ZN => n50);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n66, n67, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n100, Z => n33);
   U2 : BUF_X1 port map( A => n100, Z => n66);
   U3 : BUF_X1 port map( A => n100, Z => n67);
   U4 : INV_X1 port map( A => n101, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n33, B1 => B(0), B2 => SEL, ZN => 
                           n101);
   U6 : INV_X1 port map( A => n112, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n33, B1 => B(1), B2 => SEL, ZN => 
                           n112);
   U8 : INV_X1 port map( A => n116, ZN => Y(23));
   U9 : AOI22_X1 port map( A1 => A(23), A2 => n66, B1 => B(23), B2 => SEL, ZN 
                           => n116);
   U10 : INV_X1 port map( A => n117, ZN => Y(24));
   U11 : AOI22_X1 port map( A1 => A(24), A2 => n66, B1 => B(24), B2 => SEL, ZN 
                           => n117);
   U12 : INV_X1 port map( A => n118, ZN => Y(25));
   U13 : AOI22_X1 port map( A1 => A(25), A2 => n66, B1 => B(25), B2 => SEL, ZN 
                           => n118);
   U14 : INV_X1 port map( A => n119, ZN => Y(26));
   U15 : AOI22_X1 port map( A1 => A(26), A2 => n66, B1 => B(26), B2 => SEL, ZN 
                           => n119);
   U16 : INV_X1 port map( A => n120, ZN => Y(27));
   U17 : AOI22_X1 port map( A1 => A(27), A2 => n66, B1 => B(27), B2 => SEL, ZN 
                           => n120);
   U18 : INV_X1 port map( A => n121, ZN => Y(28));
   U19 : AOI22_X1 port map( A1 => A(28), A2 => n66, B1 => B(28), B2 => SEL, ZN 
                           => n121);
   U20 : INV_X1 port map( A => n123, ZN => Y(2));
   U21 : AOI22_X1 port map( A1 => A(2), A2 => n66, B1 => B(2), B2 => SEL, ZN =>
                           n123);
   U22 : INV_X1 port map( A => n126, ZN => Y(3));
   U23 : AOI22_X1 port map( A1 => A(3), A2 => n67, B1 => B(3), B2 => SEL, ZN =>
                           n126);
   U24 : INV_X1 port map( A => n127, ZN => Y(4));
   U25 : AOI22_X1 port map( A1 => A(4), A2 => n67, B1 => B(4), B2 => SEL, ZN =>
                           n127);
   U26 : INV_X1 port map( A => n128, ZN => Y(5));
   U27 : AOI22_X1 port map( A1 => A(5), A2 => n67, B1 => B(5), B2 => SEL, ZN =>
                           n128);
   U28 : INV_X1 port map( A => n129, ZN => Y(6));
   U29 : AOI22_X1 port map( A1 => A(6), A2 => n67, B1 => B(6), B2 => SEL, ZN =>
                           n129);
   U30 : INV_X1 port map( A => n130, ZN => Y(7));
   U31 : AOI22_X1 port map( A1 => A(7), A2 => n67, B1 => B(7), B2 => SEL, ZN =>
                           n130);
   U32 : INV_X1 port map( A => n131, ZN => Y(8));
   U33 : AOI22_X1 port map( A1 => A(8), A2 => n67, B1 => B(8), B2 => SEL, ZN =>
                           n131);
   U34 : INV_X1 port map( A => n132, ZN => Y(9));
   U35 : AOI22_X1 port map( A1 => A(9), A2 => n67, B1 => SEL, B2 => B(9), ZN =>
                           n132);
   U36 : INV_X1 port map( A => n102, ZN => Y(10));
   U37 : AOI22_X1 port map( A1 => A(10), A2 => n33, B1 => B(10), B2 => SEL, ZN 
                           => n102);
   U38 : INV_X1 port map( A => n103, ZN => Y(11));
   U39 : AOI22_X1 port map( A1 => A(11), A2 => n33, B1 => B(11), B2 => SEL, ZN 
                           => n103);
   U40 : INV_X1 port map( A => n104, ZN => Y(12));
   U41 : AOI22_X1 port map( A1 => A(12), A2 => n33, B1 => B(12), B2 => SEL, ZN 
                           => n104);
   U42 : INV_X1 port map( A => n105, ZN => Y(13));
   U43 : AOI22_X1 port map( A1 => A(13), A2 => n33, B1 => B(13), B2 => SEL, ZN 
                           => n105);
   U44 : INV_X1 port map( A => n106, ZN => Y(14));
   U45 : AOI22_X1 port map( A1 => A(14), A2 => n33, B1 => B(14), B2 => SEL, ZN 
                           => n106);
   U46 : INV_X1 port map( A => n107, ZN => Y(15));
   U47 : AOI22_X1 port map( A1 => A(15), A2 => n33, B1 => B(15), B2 => SEL, ZN 
                           => n107);
   U48 : INV_X1 port map( A => n108, ZN => Y(16));
   U49 : AOI22_X1 port map( A1 => A(16), A2 => n33, B1 => B(16), B2 => SEL, ZN 
                           => n108);
   U50 : INV_X1 port map( A => n109, ZN => Y(17));
   U51 : AOI22_X1 port map( A1 => A(17), A2 => n33, B1 => B(17), B2 => SEL, ZN 
                           => n109);
   U52 : INV_X1 port map( A => n110, ZN => Y(18));
   U53 : AOI22_X1 port map( A1 => A(18), A2 => n33, B1 => B(18), B2 => SEL, ZN 
                           => n110);
   U54 : INV_X1 port map( A => n111, ZN => Y(19));
   U55 : AOI22_X1 port map( A1 => A(19), A2 => n33, B1 => B(19), B2 => SEL, ZN 
                           => n111);
   U56 : INV_X1 port map( A => n113, ZN => Y(20));
   U57 : AOI22_X1 port map( A1 => A(20), A2 => n66, B1 => B(20), B2 => SEL, ZN 
                           => n113);
   U58 : INV_X1 port map( A => n114, ZN => Y(21));
   U59 : AOI22_X1 port map( A1 => A(21), A2 => n66, B1 => B(21), B2 => SEL, ZN 
                           => n114);
   U60 : INV_X1 port map( A => n115, ZN => Y(22));
   U61 : AOI22_X1 port map( A1 => A(22), A2 => n66, B1 => B(22), B2 => SEL, ZN 
                           => n115);
   U62 : INV_X1 port map( A => n122, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n66, B1 => B(29), B2 => SEL, ZN 
                           => n122);
   U64 : INV_X1 port map( A => n124, ZN => Y(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n66, B1 => B(30), B2 => SEL, ZN 
                           => n124);
   U66 : INV_X1 port map( A => n125, ZN => Y(31));
   U67 : AOI22_X1 port map( A1 => A(31), A2 => n67, B1 => B(31), B2 => SEL, ZN 
                           => n125);
   U68 : INV_X1 port map( A => SEL, ZN => n100);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n66, n67, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n100, Z => n33);
   U2 : BUF_X1 port map( A => n100, Z => n66);
   U3 : BUF_X1 port map( A => n100, Z => n67);
   U4 : INV_X1 port map( A => n101, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n33, B1 => B(0), B2 => SEL, ZN => 
                           n101);
   U6 : INV_X1 port map( A => n112, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n33, B1 => B(1), B2 => SEL, ZN => 
                           n112);
   U8 : INV_X1 port map( A => n116, ZN => Y(23));
   U9 : AOI22_X1 port map( A1 => A(23), A2 => n66, B1 => B(23), B2 => SEL, ZN 
                           => n116);
   U10 : INV_X1 port map( A => n117, ZN => Y(24));
   U11 : AOI22_X1 port map( A1 => A(24), A2 => n66, B1 => B(24), B2 => SEL, ZN 
                           => n117);
   U12 : INV_X1 port map( A => n118, ZN => Y(25));
   U13 : AOI22_X1 port map( A1 => A(25), A2 => n66, B1 => B(25), B2 => SEL, ZN 
                           => n118);
   U14 : INV_X1 port map( A => n119, ZN => Y(26));
   U15 : AOI22_X1 port map( A1 => A(26), A2 => n66, B1 => B(26), B2 => SEL, ZN 
                           => n119);
   U16 : INV_X1 port map( A => n120, ZN => Y(27));
   U17 : AOI22_X1 port map( A1 => A(27), A2 => n66, B1 => B(27), B2 => SEL, ZN 
                           => n120);
   U18 : INV_X1 port map( A => n121, ZN => Y(28));
   U19 : AOI22_X1 port map( A1 => A(28), A2 => n66, B1 => B(28), B2 => SEL, ZN 
                           => n121);
   U20 : INV_X1 port map( A => n123, ZN => Y(2));
   U21 : AOI22_X1 port map( A1 => A(2), A2 => n66, B1 => B(2), B2 => SEL, ZN =>
                           n123);
   U22 : INV_X1 port map( A => n126, ZN => Y(3));
   U23 : AOI22_X1 port map( A1 => A(3), A2 => n67, B1 => B(3), B2 => SEL, ZN =>
                           n126);
   U24 : INV_X1 port map( A => n127, ZN => Y(4));
   U25 : AOI22_X1 port map( A1 => A(4), A2 => n67, B1 => B(4), B2 => SEL, ZN =>
                           n127);
   U26 : INV_X1 port map( A => n128, ZN => Y(5));
   U27 : AOI22_X1 port map( A1 => A(5), A2 => n67, B1 => B(5), B2 => SEL, ZN =>
                           n128);
   U28 : INV_X1 port map( A => n129, ZN => Y(6));
   U29 : AOI22_X1 port map( A1 => A(6), A2 => n67, B1 => B(6), B2 => SEL, ZN =>
                           n129);
   U30 : INV_X1 port map( A => n130, ZN => Y(7));
   U31 : AOI22_X1 port map( A1 => A(7), A2 => n67, B1 => B(7), B2 => SEL, ZN =>
                           n130);
   U32 : INV_X1 port map( A => n131, ZN => Y(8));
   U33 : AOI22_X1 port map( A1 => A(8), A2 => n67, B1 => B(8), B2 => SEL, ZN =>
                           n131);
   U34 : INV_X1 port map( A => n132, ZN => Y(9));
   U35 : AOI22_X1 port map( A1 => A(9), A2 => n67, B1 => SEL, B2 => B(9), ZN =>
                           n132);
   U36 : INV_X1 port map( A => n102, ZN => Y(10));
   U37 : AOI22_X1 port map( A1 => A(10), A2 => n33, B1 => B(10), B2 => SEL, ZN 
                           => n102);
   U38 : INV_X1 port map( A => n103, ZN => Y(11));
   U39 : AOI22_X1 port map( A1 => A(11), A2 => n33, B1 => B(11), B2 => SEL, ZN 
                           => n103);
   U40 : INV_X1 port map( A => n104, ZN => Y(12));
   U41 : AOI22_X1 port map( A1 => A(12), A2 => n33, B1 => B(12), B2 => SEL, ZN 
                           => n104);
   U42 : INV_X1 port map( A => n105, ZN => Y(13));
   U43 : AOI22_X1 port map( A1 => A(13), A2 => n33, B1 => B(13), B2 => SEL, ZN 
                           => n105);
   U44 : INV_X1 port map( A => n106, ZN => Y(14));
   U45 : AOI22_X1 port map( A1 => A(14), A2 => n33, B1 => B(14), B2 => SEL, ZN 
                           => n106);
   U46 : INV_X1 port map( A => n107, ZN => Y(15));
   U47 : AOI22_X1 port map( A1 => A(15), A2 => n33, B1 => B(15), B2 => SEL, ZN 
                           => n107);
   U48 : INV_X1 port map( A => n108, ZN => Y(16));
   U49 : AOI22_X1 port map( A1 => A(16), A2 => n33, B1 => B(16), B2 => SEL, ZN 
                           => n108);
   U50 : INV_X1 port map( A => n109, ZN => Y(17));
   U51 : AOI22_X1 port map( A1 => A(17), A2 => n33, B1 => B(17), B2 => SEL, ZN 
                           => n109);
   U52 : INV_X1 port map( A => n110, ZN => Y(18));
   U53 : AOI22_X1 port map( A1 => A(18), A2 => n33, B1 => B(18), B2 => SEL, ZN 
                           => n110);
   U54 : INV_X1 port map( A => n111, ZN => Y(19));
   U55 : AOI22_X1 port map( A1 => A(19), A2 => n33, B1 => B(19), B2 => SEL, ZN 
                           => n111);
   U56 : INV_X1 port map( A => n113, ZN => Y(20));
   U57 : AOI22_X1 port map( A1 => A(20), A2 => n66, B1 => B(20), B2 => SEL, ZN 
                           => n113);
   U58 : INV_X1 port map( A => n114, ZN => Y(21));
   U59 : AOI22_X1 port map( A1 => A(21), A2 => n66, B1 => B(21), B2 => SEL, ZN 
                           => n114);
   U60 : INV_X1 port map( A => n115, ZN => Y(22));
   U61 : AOI22_X1 port map( A1 => A(22), A2 => n66, B1 => B(22), B2 => SEL, ZN 
                           => n115);
   U62 : INV_X1 port map( A => n122, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n66, B1 => B(29), B2 => SEL, ZN 
                           => n122);
   U64 : INV_X1 port map( A => n124, ZN => Y(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n66, B1 => B(30), B2 => SEL, ZN 
                           => n124);
   U66 : INV_X1 port map( A => n125, ZN => Y(31));
   U67 : AOI22_X1 port map( A1 => A(31), A2 => n67, B1 => B(31), B2 => SEL, ZN 
                           => n125);
   U68 : INV_X1 port map( A => SEL, ZN => n100);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n33, n66, n67, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n100, Z => n33);
   U2 : BUF_X1 port map( A => n100, Z => n66);
   U3 : BUF_X1 port map( A => n100, Z => n67);
   U4 : INV_X1 port map( A => n34, ZN => Y(9));
   U5 : AOI22_X1 port map( A1 => A(9), A2 => n67, B1 => SEL, B2 => B(9), ZN => 
                           n34);
   U6 : INV_X1 port map( A => n65, ZN => Y(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n33, B1 => B(0), B2 => SEL, ZN => 
                           n65);
   U8 : INV_X1 port map( A => n54, ZN => Y(1));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n33, B1 => B(1), B2 => SEL, ZN => 
                           n54);
   U10 : INV_X1 port map( A => n43, ZN => Y(2));
   U11 : AOI22_X1 port map( A1 => A(2), A2 => n66, B1 => B(2), B2 => SEL, ZN =>
                           n43);
   U12 : INV_X1 port map( A => n40, ZN => Y(3));
   U13 : AOI22_X1 port map( A1 => A(3), A2 => n67, B1 => B(3), B2 => SEL, ZN =>
                           n40);
   U14 : INV_X1 port map( A => n39, ZN => Y(4));
   U15 : AOI22_X1 port map( A1 => A(4), A2 => n67, B1 => B(4), B2 => SEL, ZN =>
                           n39);
   U16 : INV_X1 port map( A => n38, ZN => Y(5));
   U17 : AOI22_X1 port map( A1 => A(5), A2 => n67, B1 => B(5), B2 => SEL, ZN =>
                           n38);
   U18 : INV_X1 port map( A => n37, ZN => Y(6));
   U19 : AOI22_X1 port map( A1 => A(6), A2 => n67, B1 => B(6), B2 => SEL, ZN =>
                           n37);
   U20 : INV_X1 port map( A => n36, ZN => Y(7));
   U21 : AOI22_X1 port map( A1 => A(7), A2 => n67, B1 => B(7), B2 => SEL, ZN =>
                           n36);
   U22 : INV_X1 port map( A => n35, ZN => Y(8));
   U23 : AOI22_X1 port map( A1 => A(8), A2 => n67, B1 => B(8), B2 => SEL, ZN =>
                           n35);
   U24 : INV_X1 port map( A => n64, ZN => Y(10));
   U25 : AOI22_X1 port map( A1 => A(10), A2 => n33, B1 => B(10), B2 => SEL, ZN 
                           => n64);
   U26 : INV_X1 port map( A => n63, ZN => Y(11));
   U27 : AOI22_X1 port map( A1 => A(11), A2 => n33, B1 => B(11), B2 => SEL, ZN 
                           => n63);
   U28 : INV_X1 port map( A => n62, ZN => Y(12));
   U29 : AOI22_X1 port map( A1 => A(12), A2 => n33, B1 => B(12), B2 => SEL, ZN 
                           => n62);
   U30 : INV_X1 port map( A => n61, ZN => Y(13));
   U31 : AOI22_X1 port map( A1 => A(13), A2 => n33, B1 => B(13), B2 => SEL, ZN 
                           => n61);
   U32 : INV_X1 port map( A => n60, ZN => Y(14));
   U33 : AOI22_X1 port map( A1 => A(14), A2 => n33, B1 => B(14), B2 => SEL, ZN 
                           => n60);
   U34 : INV_X1 port map( A => n59, ZN => Y(15));
   U35 : AOI22_X1 port map( A1 => A(15), A2 => n33, B1 => B(15), B2 => SEL, ZN 
                           => n59);
   U36 : INV_X1 port map( A => n58, ZN => Y(16));
   U37 : AOI22_X1 port map( A1 => A(16), A2 => n33, B1 => B(16), B2 => SEL, ZN 
                           => n58);
   U38 : INV_X1 port map( A => n57, ZN => Y(17));
   U39 : AOI22_X1 port map( A1 => A(17), A2 => n33, B1 => B(17), B2 => SEL, ZN 
                           => n57);
   U40 : INV_X1 port map( A => n56, ZN => Y(18));
   U41 : AOI22_X1 port map( A1 => A(18), A2 => n33, B1 => B(18), B2 => SEL, ZN 
                           => n56);
   U42 : INV_X1 port map( A => n55, ZN => Y(19));
   U43 : AOI22_X1 port map( A1 => A(19), A2 => n33, B1 => B(19), B2 => SEL, ZN 
                           => n55);
   U44 : INV_X1 port map( A => n53, ZN => Y(20));
   U45 : AOI22_X1 port map( A1 => A(20), A2 => n66, B1 => B(20), B2 => SEL, ZN 
                           => n53);
   U46 : INV_X1 port map( A => n52, ZN => Y(21));
   U47 : AOI22_X1 port map( A1 => A(21), A2 => n66, B1 => B(21), B2 => SEL, ZN 
                           => n52);
   U48 : INV_X1 port map( A => n51, ZN => Y(22));
   U49 : AOI22_X1 port map( A1 => A(22), A2 => n66, B1 => B(22), B2 => SEL, ZN 
                           => n51);
   U50 : INV_X1 port map( A => n50, ZN => Y(23));
   U51 : AOI22_X1 port map( A1 => A(23), A2 => n66, B1 => B(23), B2 => SEL, ZN 
                           => n50);
   U52 : INV_X1 port map( A => n49, ZN => Y(24));
   U53 : AOI22_X1 port map( A1 => A(24), A2 => n66, B1 => B(24), B2 => SEL, ZN 
                           => n49);
   U54 : INV_X1 port map( A => n48, ZN => Y(25));
   U55 : AOI22_X1 port map( A1 => A(25), A2 => n66, B1 => B(25), B2 => SEL, ZN 
                           => n48);
   U56 : INV_X1 port map( A => n47, ZN => Y(26));
   U57 : AOI22_X1 port map( A1 => A(26), A2 => n66, B1 => B(26), B2 => SEL, ZN 
                           => n47);
   U58 : INV_X1 port map( A => n46, ZN => Y(27));
   U59 : AOI22_X1 port map( A1 => A(27), A2 => n66, B1 => B(27), B2 => SEL, ZN 
                           => n46);
   U60 : INV_X1 port map( A => n45, ZN => Y(28));
   U61 : AOI22_X1 port map( A1 => A(28), A2 => n66, B1 => B(28), B2 => SEL, ZN 
                           => n45);
   U62 : INV_X1 port map( A => n44, ZN => Y(29));
   U63 : AOI22_X1 port map( A1 => A(29), A2 => n66, B1 => B(29), B2 => SEL, ZN 
                           => n44);
   U64 : INV_X1 port map( A => n42, ZN => Y(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n66, B1 => B(30), B2 => SEL, ZN 
                           => n42);
   U66 : INV_X1 port map( A => n41, ZN => Y(31));
   U67 : AOI22_X1 port map( A1 => A(31), A2 => n67, B1 => B(31), B2 => SEL, ZN 
                           => n41);
   U68 : INV_X1 port map( A => SEL, ZN => n100);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity branch_block_nbit32 is

   port( branch_op : in std_logic;  cmp_out, PC, label_PC : in std_logic_vector
         (31 downto 0);  next_PC : out std_logic_vector (31 downto 0));

end branch_block_nbit32;

architecture SYN_struct of branch_block_nbit32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal branch_taken : std_logic;

begin
   
   next_pc_mux : MUX21_GENERIC_NBIT32_1 port map( A(31) => PC(31), A(30) => 
                           PC(30), A(29) => PC(29), A(28) => PC(28), A(27) => 
                           PC(27), A(26) => PC(26), A(25) => PC(25), A(24) => 
                           PC(24), A(23) => PC(23), A(22) => PC(22), A(21) => 
                           PC(21), A(20) => PC(20), A(19) => PC(19), A(18) => 
                           PC(18), A(17) => PC(17), A(16) => PC(16), A(15) => 
                           PC(15), A(14) => PC(14), A(13) => PC(13), A(12) => 
                           PC(12), A(11) => PC(11), A(10) => PC(10), A(9) => 
                           PC(9), A(8) => PC(8), A(7) => PC(7), A(6) => PC(6), 
                           A(5) => PC(5), A(4) => PC(4), A(3) => PC(3), A(2) =>
                           PC(2), A(1) => PC(1), A(0) => PC(0), B(31) => 
                           label_PC(31), B(30) => label_PC(30), B(29) => 
                           label_PC(29), B(28) => label_PC(28), B(27) => 
                           label_PC(27), B(26) => label_PC(26), B(25) => 
                           label_PC(25), B(24) => label_PC(24), B(23) => 
                           label_PC(23), B(22) => label_PC(22), B(21) => 
                           label_PC(21), B(20) => label_PC(20), B(19) => 
                           label_PC(19), B(18) => label_PC(18), B(17) => 
                           label_PC(17), B(16) => label_PC(16), B(15) => 
                           label_PC(15), B(14) => label_PC(14), B(13) => 
                           label_PC(13), B(12) => label_PC(12), B(11) => 
                           label_PC(11), B(10) => label_PC(10), B(9) => 
                           label_PC(9), B(8) => label_PC(8), B(7) => 
                           label_PC(7), B(6) => label_PC(6), B(5) => 
                           label_PC(5), B(4) => label_PC(4), B(3) => 
                           label_PC(3), B(2) => label_PC(2), B(1) => 
                           label_PC(1), B(0) => label_PC(0), SEL => 
                           branch_taken, Y(31) => next_PC(31), Y(30) => 
                           next_PC(30), Y(29) => next_PC(29), Y(28) => 
                           next_PC(28), Y(27) => next_PC(27), Y(26) => 
                           next_PC(26), Y(25) => next_PC(25), Y(24) => 
                           next_PC(24), Y(23) => next_PC(23), Y(22) => 
                           next_PC(22), Y(21) => next_PC(21), Y(20) => 
                           next_PC(20), Y(19) => next_PC(19), Y(18) => 
                           next_PC(18), Y(17) => next_PC(17), Y(16) => 
                           next_PC(16), Y(15) => next_PC(15), Y(14) => 
                           next_PC(14), Y(13) => next_PC(13), Y(12) => 
                           next_PC(12), Y(11) => next_PC(11), Y(10) => 
                           next_PC(10), Y(9) => next_PC(9), Y(8) => next_PC(8),
                           Y(7) => next_PC(7), Y(6) => next_PC(6), Y(5) => 
                           next_PC(5), Y(4) => next_PC(4), Y(3) => next_PC(3), 
                           Y(2) => next_PC(2), Y(1) => next_PC(1), Y(0) => 
                           next_PC(0));
   U1 : AND2_X1 port map( A1 => cmp_out(0), A2 => branch_op, ZN => branch_taken
                           );

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_4 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_4;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n52, Q => Q(31), 
                           QN => n148);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n52, Q => Q(30), 
                           QN => n147);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n52, Q => Q(29), 
                           QN => n146);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n52, Q => Q(28), 
                           QN => n145);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n52, Q => Q(27), 
                           QN => n144);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n52, Q => Q(26), 
                           QN => n143);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n52, Q => Q(25),
                           QN => n142);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n52, Q => Q(24),
                           QN => n141);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n51, Q => Q(23),
                           QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n51, Q => Q(22),
                           QN => n139);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n51, Q => Q(21),
                           QN => n138);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n51, Q => Q(20),
                           QN => n137);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n136);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n135);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n51, Q => Q(17),
                           QN => n134);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n133);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n132);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n131);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n51, Q => Q(13),
                           QN => n130);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n51, Q => Q(12),
                           QN => n129);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n50, Q => Q(11),
                           QN => n128);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n50, Q => Q(10),
                           QN => n127);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n50, Q => Q(9), 
                           QN => n126);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n50, Q => Q(8), 
                           QN => n125);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n50, Q => Q(7), 
                           QN => n124);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n50, Q => Q(6), 
                           QN => n123);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n50, Q => Q(5), 
                           QN => n122);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n50, Q => Q(4), 
                           QN => n121);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n50, Q => Q(3), 
                           QN => n120);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n50, Q => Q(2), 
                           QN => n119);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n50, Q => Q(1), 
                           QN => n118);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n50, Q => Q(0), 
                           QN => n117);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n50);
   U5 : BUF_X1 port map( A => RESET_n, Z => n51);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n44);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n117, A2 => n40, B1 => n42, B2 => n116, ZN =>
                           n35);
   U20 : INV_X1 port map( A => D(0), ZN => n116);
   U21 : OAI22_X1 port map( A1 => n118, A2 => n39, B1 => n42, B2 => n115, ZN =>
                           n34);
   U22 : INV_X1 port map( A => D(1), ZN => n115);
   U23 : OAI22_X1 port map( A1 => n143, A2 => n40, B1 => n41, B2 => n58, ZN => 
                           n9);
   U24 : INV_X1 port map( A => D(26), ZN => n58);
   U25 : OAI22_X1 port map( A1 => n144, A2 => n39, B1 => n41, B2 => n57, ZN => 
                           n8);
   U26 : INV_X1 port map( A => D(27), ZN => n57);
   U27 : OAI22_X1 port map( A1 => n145, A2 => n40, B1 => n41, B2 => n56, ZN => 
                           n7);
   U28 : INV_X1 port map( A => D(28), ZN => n56);
   U29 : OAI22_X1 port map( A1 => n146, A2 => n39, B1 => n41, B2 => n55, ZN => 
                           n6);
   U30 : INV_X1 port map( A => D(29), ZN => n55);
   U31 : OAI22_X1 port map( A1 => n147, A2 => n40, B1 => n42, B2 => n54, ZN => 
                           n5);
   U32 : INV_X1 port map( A => D(30), ZN => n54);
   U33 : OAI22_X1 port map( A1 => n148, A2 => n39, B1 => n42, B2 => n53, ZN => 
                           n4);
   U34 : INV_X1 port map( A => D(31), ZN => n53);
   U35 : OAI22_X1 port map( A1 => n129, A2 => n40, B1 => n45, B2 => n104, ZN =>
                           n23);
   U36 : INV_X1 port map( A => D(12), ZN => n104);
   U37 : OAI22_X1 port map( A1 => n130, A2 => n40, B1 => n45, B2 => n103, ZN =>
                           n22);
   U38 : INV_X1 port map( A => D(13), ZN => n103);
   U39 : OAI22_X1 port map( A1 => n131, A2 => n39, B1 => n46, B2 => n102, ZN =>
                           n21);
   U40 : INV_X1 port map( A => D(14), ZN => n102);
   U41 : OAI22_X1 port map( A1 => n132, A2 => n39, B1 => n46, B2 => n101, ZN =>
                           n20);
   U42 : INV_X1 port map( A => D(15), ZN => n101);
   U43 : OAI22_X1 port map( A1 => n133, A2 => n39, B1 => n46, B2 => n100, ZN =>
                           n19);
   U44 : INV_X1 port map( A => D(16), ZN => n100);
   U45 : OAI22_X1 port map( A1 => n134, A2 => n39, B1 => n46, B2 => n99, ZN => 
                           n18);
   U46 : INV_X1 port map( A => D(17), ZN => n99);
   U47 : OAI22_X1 port map( A1 => n135, A2 => n39, B1 => n47, B2 => n98, ZN => 
                           n17);
   U48 : INV_X1 port map( A => D(18), ZN => n98);
   U49 : OAI22_X1 port map( A1 => n136, A2 => n39, B1 => n47, B2 => n65, ZN => 
                           n16);
   U50 : INV_X1 port map( A => D(19), ZN => n65);
   U51 : OAI22_X1 port map( A1 => n137, A2 => n39, B1 => n47, B2 => n64, ZN => 
                           n15);
   U52 : INV_X1 port map( A => D(20), ZN => n64);
   U53 : OAI22_X1 port map( A1 => n138, A2 => n39, B1 => n47, B2 => n63, ZN => 
                           n14);
   U54 : INV_X1 port map( A => D(21), ZN => n63);
   U55 : OAI22_X1 port map( A1 => n139, A2 => n39, B1 => n48, B2 => n62, ZN => 
                           n13);
   U56 : INV_X1 port map( A => D(22), ZN => n62);
   U57 : OAI22_X1 port map( A1 => n140, A2 => n39, B1 => n48, B2 => n61, ZN => 
                           n12);
   U58 : INV_X1 port map( A => D(23), ZN => n61);
   U59 : OAI22_X1 port map( A1 => n141, A2 => n39, B1 => n48, B2 => n60, ZN => 
                           n11);
   U60 : INV_X1 port map( A => D(24), ZN => n60);
   U61 : OAI22_X1 port map( A1 => n142, A2 => n39, B1 => n48, B2 => n59, ZN => 
                           n10);
   U62 : INV_X1 port map( A => D(25), ZN => n59);
   U63 : OAI22_X1 port map( A1 => n119, A2 => n40, B1 => n43, B2 => n114, ZN =>
                           n33);
   U64 : INV_X1 port map( A => D(2), ZN => n114);
   U65 : OAI22_X1 port map( A1 => n120, A2 => n40, B1 => n43, B2 => n113, ZN =>
                           n32);
   U66 : INV_X1 port map( A => D(3), ZN => n113);
   U67 : OAI22_X1 port map( A1 => n121, A2 => n40, B1 => n43, B2 => n112, ZN =>
                           n31);
   U68 : INV_X1 port map( A => D(4), ZN => n112);
   U69 : OAI22_X1 port map( A1 => n122, A2 => n40, B1 => n43, B2 => n111, ZN =>
                           n30);
   U70 : INV_X1 port map( A => D(5), ZN => n111);
   U71 : OAI22_X1 port map( A1 => n123, A2 => n40, B1 => n44, B2 => n110, ZN =>
                           n29);
   U72 : INV_X1 port map( A => D(6), ZN => n110);
   U73 : OAI22_X1 port map( A1 => n124, A2 => n40, B1 => n44, B2 => n109, ZN =>
                           n28);
   U74 : INV_X1 port map( A => D(7), ZN => n109);
   U75 : OAI22_X1 port map( A1 => n125, A2 => n40, B1 => n44, B2 => n108, ZN =>
                           n27);
   U76 : INV_X1 port map( A => D(8), ZN => n108);
   U77 : OAI22_X1 port map( A1 => n126, A2 => n40, B1 => n44, B2 => n107, ZN =>
                           n26);
   U78 : INV_X1 port map( A => D(9), ZN => n107);
   U79 : OAI22_X1 port map( A1 => n127, A2 => n40, B1 => n45, B2 => n106, ZN =>
                           n25);
   U80 : INV_X1 port map( A => D(10), ZN => n106);
   U81 : OAI22_X1 port map( A1 => n128, A2 => n40, B1 => n45, B2 => n105, ZN =>
                           n24);
   U82 : INV_X1 port map( A => D(11), ZN => n105);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_5 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_5;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n50, Q => Q(31), 
                           QN => n148);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n50, Q => Q(30), 
                           QN => n147);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n50, Q => Q(29), 
                           QN => n146);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n50, Q => Q(28), 
                           QN => n145);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n50, Q => Q(27), 
                           QN => n144);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n50, Q => Q(26), 
                           QN => n143);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n50, Q => Q(25),
                           QN => n142);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n50, Q => Q(24),
                           QN => n141);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n50, Q => Q(23),
                           QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n50, Q => Q(22),
                           QN => n139);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n50, Q => Q(21),
                           QN => n138);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n50, Q => Q(20),
                           QN => n137);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n136);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n135);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n51, Q => Q(17),
                           QN => n134);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n133);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n132);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n131);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n51, Q => Q(13),
                           QN => n130);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n51, Q => Q(12),
                           QN => n129);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n51, Q => Q(11),
                           QN => n128);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n51, Q => Q(10),
                           QN => n127);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n51, Q => Q(9), 
                           QN => n126);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n51, Q => Q(8), 
                           QN => n125);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n52, Q => Q(7), 
                           QN => n124);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n52, Q => Q(6), 
                           QN => n123);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n52, Q => Q(5), 
                           QN => n122);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n52, Q => Q(4), 
                           QN => n121);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n52, Q => Q(3), 
                           QN => n120);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n52, Q => Q(2), 
                           QN => n119);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n52, Q => Q(1), 
                           QN => n118);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n52, Q => Q(0), 
                           QN => n117);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n51);
   U5 : BUF_X1 port map( A => RESET_n, Z => n50);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n44);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n117, A2 => n40, B1 => n42, B2 => n116, ZN =>
                           n35);
   U20 : INV_X1 port map( A => D(0), ZN => n116);
   U21 : OAI22_X1 port map( A1 => n118, A2 => n39, B1 => n42, B2 => n115, ZN =>
                           n34);
   U22 : INV_X1 port map( A => D(1), ZN => n115);
   U23 : OAI22_X1 port map( A1 => n143, A2 => n40, B1 => n41, B2 => n58, ZN => 
                           n9);
   U24 : INV_X1 port map( A => D(26), ZN => n58);
   U25 : OAI22_X1 port map( A1 => n144, A2 => n39, B1 => n41, B2 => n57, ZN => 
                           n8);
   U26 : INV_X1 port map( A => D(27), ZN => n57);
   U27 : OAI22_X1 port map( A1 => n145, A2 => n40, B1 => n41, B2 => n56, ZN => 
                           n7);
   U28 : INV_X1 port map( A => D(28), ZN => n56);
   U29 : OAI22_X1 port map( A1 => n146, A2 => n39, B1 => n41, B2 => n55, ZN => 
                           n6);
   U30 : INV_X1 port map( A => D(29), ZN => n55);
   U31 : OAI22_X1 port map( A1 => n147, A2 => n40, B1 => n42, B2 => n54, ZN => 
                           n5);
   U32 : INV_X1 port map( A => D(30), ZN => n54);
   U33 : OAI22_X1 port map( A1 => n148, A2 => n39, B1 => n42, B2 => n53, ZN => 
                           n4);
   U34 : INV_X1 port map( A => D(31), ZN => n53);
   U35 : OAI22_X1 port map( A1 => n119, A2 => n40, B1 => n43, B2 => n114, ZN =>
                           n33);
   U36 : INV_X1 port map( A => D(2), ZN => n114);
   U37 : OAI22_X1 port map( A1 => n120, A2 => n40, B1 => n43, B2 => n113, ZN =>
                           n32);
   U38 : INV_X1 port map( A => D(3), ZN => n113);
   U39 : OAI22_X1 port map( A1 => n121, A2 => n40, B1 => n43, B2 => n112, ZN =>
                           n31);
   U40 : INV_X1 port map( A => D(4), ZN => n112);
   U41 : OAI22_X1 port map( A1 => n122, A2 => n40, B1 => n43, B2 => n111, ZN =>
                           n30);
   U42 : INV_X1 port map( A => D(5), ZN => n111);
   U43 : OAI22_X1 port map( A1 => n123, A2 => n40, B1 => n44, B2 => n110, ZN =>
                           n29);
   U44 : INV_X1 port map( A => D(6), ZN => n110);
   U45 : OAI22_X1 port map( A1 => n124, A2 => n40, B1 => n44, B2 => n109, ZN =>
                           n28);
   U46 : INV_X1 port map( A => D(7), ZN => n109);
   U47 : OAI22_X1 port map( A1 => n125, A2 => n40, B1 => n44, B2 => n108, ZN =>
                           n27);
   U48 : INV_X1 port map( A => D(8), ZN => n108);
   U49 : OAI22_X1 port map( A1 => n126, A2 => n40, B1 => n44, B2 => n107, ZN =>
                           n26);
   U50 : INV_X1 port map( A => D(9), ZN => n107);
   U51 : OAI22_X1 port map( A1 => n127, A2 => n40, B1 => n45, B2 => n106, ZN =>
                           n25);
   U52 : INV_X1 port map( A => D(10), ZN => n106);
   U53 : OAI22_X1 port map( A1 => n128, A2 => n40, B1 => n45, B2 => n105, ZN =>
                           n24);
   U54 : INV_X1 port map( A => D(11), ZN => n105);
   U55 : OAI22_X1 port map( A1 => n129, A2 => n40, B1 => n45, B2 => n104, ZN =>
                           n23);
   U56 : INV_X1 port map( A => D(12), ZN => n104);
   U57 : OAI22_X1 port map( A1 => n130, A2 => n40, B1 => n45, B2 => n103, ZN =>
                           n22);
   U58 : INV_X1 port map( A => D(13), ZN => n103);
   U59 : OAI22_X1 port map( A1 => n131, A2 => n39, B1 => n46, B2 => n102, ZN =>
                           n21);
   U60 : INV_X1 port map( A => D(14), ZN => n102);
   U61 : OAI22_X1 port map( A1 => n132, A2 => n39, B1 => n46, B2 => n101, ZN =>
                           n20);
   U62 : INV_X1 port map( A => D(15), ZN => n101);
   U63 : OAI22_X1 port map( A1 => n133, A2 => n39, B1 => n46, B2 => n100, ZN =>
                           n19);
   U64 : INV_X1 port map( A => D(16), ZN => n100);
   U65 : OAI22_X1 port map( A1 => n134, A2 => n39, B1 => n46, B2 => n99, ZN => 
                           n18);
   U66 : INV_X1 port map( A => D(17), ZN => n99);
   U67 : OAI22_X1 port map( A1 => n135, A2 => n39, B1 => n47, B2 => n98, ZN => 
                           n17);
   U68 : INV_X1 port map( A => D(18), ZN => n98);
   U69 : OAI22_X1 port map( A1 => n136, A2 => n39, B1 => n47, B2 => n65, ZN => 
                           n16);
   U70 : INV_X1 port map( A => D(19), ZN => n65);
   U71 : OAI22_X1 port map( A1 => n137, A2 => n39, B1 => n47, B2 => n64, ZN => 
                           n15);
   U72 : INV_X1 port map( A => D(20), ZN => n64);
   U73 : OAI22_X1 port map( A1 => n138, A2 => n39, B1 => n47, B2 => n63, ZN => 
                           n14);
   U74 : INV_X1 port map( A => D(21), ZN => n63);
   U75 : OAI22_X1 port map( A1 => n139, A2 => n39, B1 => n48, B2 => n62, ZN => 
                           n13);
   U76 : INV_X1 port map( A => D(22), ZN => n62);
   U77 : OAI22_X1 port map( A1 => n140, A2 => n39, B1 => n48, B2 => n61, ZN => 
                           n12);
   U78 : INV_X1 port map( A => D(23), ZN => n61);
   U79 : OAI22_X1 port map( A1 => n141, A2 => n39, B1 => n48, B2 => n60, ZN => 
                           n11);
   U80 : INV_X1 port map( A => D(24), ZN => n60);
   U81 : OAI22_X1 port map( A1 => n142, A2 => n39, B1 => n48, B2 => n59, ZN => 
                           n10);
   U82 : INV_X1 port map( A => D(25), ZN => n59);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_6 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_6;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n50, Q => Q(31), 
                           QN => n148);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n50, Q => Q(30), 
                           QN => n147);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n50, Q => Q(29), 
                           QN => n146);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n50, Q => Q(28), 
                           QN => n145);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n50, Q => Q(27), 
                           QN => n144);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n50, Q => Q(26), 
                           QN => n143);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n50, Q => Q(25),
                           QN => n142);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n50, Q => Q(24),
                           QN => n141);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n50, Q => Q(23),
                           QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n50, Q => Q(22),
                           QN => n139);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n50, Q => Q(21),
                           QN => n138);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n50, Q => Q(20),
                           QN => n137);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n136);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n135);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n51, Q => Q(17),
                           QN => n134);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n133);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n132);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n131);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n51, Q => Q(13),
                           QN => n130);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n51, Q => Q(12),
                           QN => n129);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n51, Q => Q(11),
                           QN => n128);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n51, Q => Q(10),
                           QN => n127);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n51, Q => Q(9), 
                           QN => n126);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n51, Q => Q(8), 
                           QN => n125);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n52, Q => Q(7), 
                           QN => n124);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n52, Q => Q(6), 
                           QN => n123);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n52, Q => Q(5), 
                           QN => n122);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n52, Q => Q(4), 
                           QN => n121);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n52, Q => Q(3), 
                           QN => n120);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n52, Q => Q(2), 
                           QN => n119);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n52, Q => Q(1), 
                           QN => n118);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n52, Q => Q(0), 
                           QN => n117);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n51);
   U5 : BUF_X1 port map( A => RESET_n, Z => n50);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n44);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n136, A2 => n39, B1 => n47, B2 => n101, ZN =>
                           n16);
   U20 : INV_X1 port map( A => D(19), ZN => n101);
   U21 : OAI22_X1 port map( A1 => n129, A2 => n40, B1 => n45, B2 => n100, ZN =>
                           n23);
   U22 : INV_X1 port map( A => D(12), ZN => n100);
   U23 : OAI22_X1 port map( A1 => n130, A2 => n40, B1 => n45, B2 => n99, ZN => 
                           n22);
   U24 : INV_X1 port map( A => D(13), ZN => n99);
   U25 : OAI22_X1 port map( A1 => n131, A2 => n39, B1 => n46, B2 => n98, ZN => 
                           n21);
   U26 : INV_X1 port map( A => D(14), ZN => n98);
   U27 : OAI22_X1 port map( A1 => n132, A2 => n39, B1 => n46, B2 => n65, ZN => 
                           n20);
   U28 : INV_X1 port map( A => D(15), ZN => n65);
   U29 : OAI22_X1 port map( A1 => n137, A2 => n39, B1 => n47, B2 => n108, ZN =>
                           n15);
   U30 : INV_X1 port map( A => D(20), ZN => n108);
   U31 : OAI22_X1 port map( A1 => n138, A2 => n39, B1 => n47, B2 => n107, ZN =>
                           n14);
   U32 : INV_X1 port map( A => D(21), ZN => n107);
   U33 : OAI22_X1 port map( A1 => n139, A2 => n39, B1 => n48, B2 => n106, ZN =>
                           n13);
   U34 : INV_X1 port map( A => D(22), ZN => n106);
   U35 : OAI22_X1 port map( A1 => n140, A2 => n39, B1 => n48, B2 => n105, ZN =>
                           n12);
   U36 : INV_X1 port map( A => D(23), ZN => n105);
   U37 : OAI22_X1 port map( A1 => n141, A2 => n39, B1 => n48, B2 => n112, ZN =>
                           n11);
   U38 : INV_X1 port map( A => D(24), ZN => n112);
   U39 : OAI22_X1 port map( A1 => n142, A2 => n39, B1 => n48, B2 => n111, ZN =>
                           n10);
   U40 : INV_X1 port map( A => D(25), ZN => n111);
   U41 : OAI22_X1 port map( A1 => n143, A2 => n40, B1 => n41, B2 => n110, ZN =>
                           n9);
   U42 : INV_X1 port map( A => D(26), ZN => n110);
   U43 : OAI22_X1 port map( A1 => n144, A2 => n39, B1 => n41, B2 => n109, ZN =>
                           n8);
   U44 : INV_X1 port map( A => D(27), ZN => n109);
   U45 : OAI22_X1 port map( A1 => n145, A2 => n40, B1 => n41, B2 => n116, ZN =>
                           n7);
   U46 : INV_X1 port map( A => D(28), ZN => n116);
   U47 : OAI22_X1 port map( A1 => n146, A2 => n39, B1 => n41, B2 => n115, ZN =>
                           n6);
   U48 : INV_X1 port map( A => D(29), ZN => n115);
   U49 : OAI22_X1 port map( A1 => n147, A2 => n40, B1 => n42, B2 => n114, ZN =>
                           n5);
   U50 : INV_X1 port map( A => D(30), ZN => n114);
   U51 : OAI22_X1 port map( A1 => n148, A2 => n39, B1 => n42, B2 => n113, ZN =>
                           n4);
   U52 : INV_X1 port map( A => D(31), ZN => n113);
   U53 : OAI22_X1 port map( A1 => n133, A2 => n39, B1 => n46, B2 => n104, ZN =>
                           n19);
   U54 : INV_X1 port map( A => D(16), ZN => n104);
   U55 : OAI22_X1 port map( A1 => n134, A2 => n39, B1 => n46, B2 => n103, ZN =>
                           n18);
   U56 : INV_X1 port map( A => D(17), ZN => n103);
   U57 : OAI22_X1 port map( A1 => n135, A2 => n39, B1 => n47, B2 => n102, ZN =>
                           n17);
   U58 : INV_X1 port map( A => D(18), ZN => n102);
   U59 : OAI22_X1 port map( A1 => n117, A2 => n40, B1 => n42, B2 => n56, ZN => 
                           n35);
   U60 : INV_X1 port map( A => D(0), ZN => n56);
   U61 : OAI22_X1 port map( A1 => n125, A2 => n40, B1 => n44, B2 => n64, ZN => 
                           n27);
   U62 : INV_X1 port map( A => D(8), ZN => n64);
   U63 : OAI22_X1 port map( A1 => n126, A2 => n40, B1 => n44, B2 => n63, ZN => 
                           n26);
   U64 : INV_X1 port map( A => D(9), ZN => n63);
   U65 : OAI22_X1 port map( A1 => n127, A2 => n40, B1 => n45, B2 => n62, ZN => 
                           n25);
   U66 : INV_X1 port map( A => D(10), ZN => n62);
   U67 : OAI22_X1 port map( A1 => n121, A2 => n40, B1 => n43, B2 => n60, ZN => 
                           n31);
   U68 : INV_X1 port map( A => D(4), ZN => n60);
   U69 : OAI22_X1 port map( A1 => n122, A2 => n40, B1 => n43, B2 => n59, ZN => 
                           n30);
   U70 : INV_X1 port map( A => D(5), ZN => n59);
   U71 : OAI22_X1 port map( A1 => n123, A2 => n40, B1 => n44, B2 => n58, ZN => 
                           n29);
   U72 : INV_X1 port map( A => D(6), ZN => n58);
   U73 : OAI22_X1 port map( A1 => n128, A2 => n40, B1 => n45, B2 => n61, ZN => 
                           n24);
   U74 : INV_X1 port map( A => D(11), ZN => n61);
   U75 : OAI22_X1 port map( A1 => n124, A2 => n40, B1 => n44, B2 => n57, ZN => 
                           n28);
   U76 : INV_X1 port map( A => D(7), ZN => n57);
   U77 : OAI22_X1 port map( A1 => n118, A2 => n39, B1 => n42, B2 => n55, ZN => 
                           n34);
   U78 : INV_X1 port map( A => D(1), ZN => n55);
   U79 : OAI22_X1 port map( A1 => n119, A2 => n40, B1 => n43, B2 => n54, ZN => 
                           n33);
   U80 : INV_X1 port map( A => D(2), ZN => n54);
   U81 : OAI22_X1 port map( A1 => n120, A2 => n40, B1 => n43, B2 => n53, ZN => 
                           n32);
   U82 : INV_X1 port map( A => D(3), ZN => n53);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_7 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_7;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n50, Q => Q(31), 
                           QN => n148);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n50, Q => Q(30), 
                           QN => n147);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n50, Q => Q(29), 
                           QN => n146);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n50, Q => Q(28), 
                           QN => n145);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n50, Q => Q(27), 
                           QN => n144);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n50, Q => Q(26), 
                           QN => n143);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n50, Q => Q(25),
                           QN => n142);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n50, Q => Q(24),
                           QN => n141);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n50, Q => Q(23),
                           QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n50, Q => Q(22),
                           QN => n139);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n50, Q => Q(21),
                           QN => n138);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n50, Q => Q(20),
                           QN => n137);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n136);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n135);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n51, Q => Q(17),
                           QN => n134);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n133);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n132);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n131);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n51, Q => Q(13),
                           QN => n130);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n51, Q => Q(12),
                           QN => n129);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n51, Q => Q(11),
                           QN => n128);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n51, Q => Q(10),
                           QN => n127);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n51, Q => Q(9), 
                           QN => n126);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n51, Q => Q(8), 
                           QN => n125);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n52, Q => Q(7), 
                           QN => n124);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n52, Q => Q(6), 
                           QN => n123);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n52, Q => Q(5), 
                           QN => n122);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n52, Q => Q(4), 
                           QN => n121);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n52, Q => Q(3), 
                           QN => n120);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n52, Q => Q(2), 
                           QN => n119);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n52, Q => Q(1), 
                           QN => n118);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n52, Q => Q(0), 
                           QN => n117);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n51);
   U5 : BUF_X1 port map( A => RESET_n, Z => n50);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n44);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n136, A2 => n39, B1 => n47, B2 => n101, ZN =>
                           n16);
   U20 : INV_X1 port map( A => D(19), ZN => n101);
   U21 : OAI22_X1 port map( A1 => n129, A2 => n40, B1 => n45, B2 => n100, ZN =>
                           n23);
   U22 : INV_X1 port map( A => D(12), ZN => n100);
   U23 : OAI22_X1 port map( A1 => n130, A2 => n40, B1 => n45, B2 => n99, ZN => 
                           n22);
   U24 : INV_X1 port map( A => D(13), ZN => n99);
   U25 : OAI22_X1 port map( A1 => n131, A2 => n39, B1 => n46, B2 => n98, ZN => 
                           n21);
   U26 : INV_X1 port map( A => D(14), ZN => n98);
   U27 : OAI22_X1 port map( A1 => n143, A2 => n40, B1 => n41, B2 => n110, ZN =>
                           n9);
   U28 : INV_X1 port map( A => D(26), ZN => n110);
   U29 : OAI22_X1 port map( A1 => n144, A2 => n39, B1 => n41, B2 => n109, ZN =>
                           n8);
   U30 : INV_X1 port map( A => D(27), ZN => n109);
   U31 : OAI22_X1 port map( A1 => n145, A2 => n40, B1 => n41, B2 => n116, ZN =>
                           n7);
   U32 : INV_X1 port map( A => D(28), ZN => n116);
   U33 : OAI22_X1 port map( A1 => n146, A2 => n39, B1 => n41, B2 => n115, ZN =>
                           n6);
   U34 : INV_X1 port map( A => D(29), ZN => n115);
   U35 : OAI22_X1 port map( A1 => n147, A2 => n40, B1 => n42, B2 => n114, ZN =>
                           n5);
   U36 : INV_X1 port map( A => D(30), ZN => n114);
   U37 : OAI22_X1 port map( A1 => n148, A2 => n39, B1 => n42, B2 => n113, ZN =>
                           n4);
   U38 : INV_X1 port map( A => D(31), ZN => n113);
   U39 : OAI22_X1 port map( A1 => n132, A2 => n39, B1 => n46, B2 => n65, ZN => 
                           n20);
   U40 : INV_X1 port map( A => D(15), ZN => n65);
   U41 : OAI22_X1 port map( A1 => n133, A2 => n39, B1 => n46, B2 => n104, ZN =>
                           n19);
   U42 : INV_X1 port map( A => D(16), ZN => n104);
   U43 : OAI22_X1 port map( A1 => n134, A2 => n39, B1 => n46, B2 => n103, ZN =>
                           n18);
   U44 : INV_X1 port map( A => D(17), ZN => n103);
   U45 : OAI22_X1 port map( A1 => n135, A2 => n39, B1 => n47, B2 => n102, ZN =>
                           n17);
   U46 : INV_X1 port map( A => D(18), ZN => n102);
   U47 : OAI22_X1 port map( A1 => n137, A2 => n39, B1 => n47, B2 => n108, ZN =>
                           n15);
   U48 : INV_X1 port map( A => D(20), ZN => n108);
   U49 : OAI22_X1 port map( A1 => n138, A2 => n39, B1 => n47, B2 => n107, ZN =>
                           n14);
   U50 : INV_X1 port map( A => D(21), ZN => n107);
   U51 : OAI22_X1 port map( A1 => n139, A2 => n39, B1 => n48, B2 => n106, ZN =>
                           n13);
   U52 : INV_X1 port map( A => D(22), ZN => n106);
   U53 : OAI22_X1 port map( A1 => n140, A2 => n39, B1 => n48, B2 => n105, ZN =>
                           n12);
   U54 : INV_X1 port map( A => D(23), ZN => n105);
   U55 : OAI22_X1 port map( A1 => n141, A2 => n39, B1 => n48, B2 => n112, ZN =>
                           n11);
   U56 : INV_X1 port map( A => D(24), ZN => n112);
   U57 : OAI22_X1 port map( A1 => n142, A2 => n39, B1 => n48, B2 => n111, ZN =>
                           n10);
   U58 : INV_X1 port map( A => D(25), ZN => n111);
   U59 : OAI22_X1 port map( A1 => n117, A2 => n40, B1 => n42, B2 => n56, ZN => 
                           n35);
   U60 : INV_X1 port map( A => D(0), ZN => n56);
   U61 : OAI22_X1 port map( A1 => n125, A2 => n40, B1 => n44, B2 => n64, ZN => 
                           n27);
   U62 : INV_X1 port map( A => D(8), ZN => n64);
   U63 : OAI22_X1 port map( A1 => n126, A2 => n40, B1 => n44, B2 => n63, ZN => 
                           n26);
   U64 : INV_X1 port map( A => D(9), ZN => n63);
   U65 : OAI22_X1 port map( A1 => n127, A2 => n40, B1 => n45, B2 => n62, ZN => 
                           n25);
   U66 : INV_X1 port map( A => D(10), ZN => n62);
   U67 : OAI22_X1 port map( A1 => n121, A2 => n40, B1 => n43, B2 => n60, ZN => 
                           n31);
   U68 : INV_X1 port map( A => D(4), ZN => n60);
   U69 : OAI22_X1 port map( A1 => n122, A2 => n40, B1 => n43, B2 => n59, ZN => 
                           n30);
   U70 : INV_X1 port map( A => D(5), ZN => n59);
   U71 : OAI22_X1 port map( A1 => n123, A2 => n40, B1 => n44, B2 => n58, ZN => 
                           n29);
   U72 : INV_X1 port map( A => D(6), ZN => n58);
   U73 : OAI22_X1 port map( A1 => n128, A2 => n40, B1 => n45, B2 => n61, ZN => 
                           n24);
   U74 : INV_X1 port map( A => D(11), ZN => n61);
   U75 : OAI22_X1 port map( A1 => n124, A2 => n40, B1 => n44, B2 => n57, ZN => 
                           n28);
   U76 : INV_X1 port map( A => D(7), ZN => n57);
   U77 : OAI22_X1 port map( A1 => n118, A2 => n39, B1 => n42, B2 => n55, ZN => 
                           n34);
   U78 : INV_X1 port map( A => D(1), ZN => n55);
   U79 : OAI22_X1 port map( A1 => n119, A2 => n40, B1 => n43, B2 => n54, ZN => 
                           n33);
   U80 : INV_X1 port map( A => D(2), ZN => n54);
   U81 : OAI22_X1 port map( A1 => n120, A2 => n40, B1 => n43, B2 => n53, ZN => 
                           n32);
   U82 : INV_X1 port map( A => D(3), ZN => n53);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity P4_ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic;  Y : out std_logic_vector (31 downto 0));

end P4_ADDER_NBIT32_NBIT_PER_BLOCK4_2;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32_NBIT_PER_BLOCK4_2 is

   component SUMGEN_NBIT32_NBLOCKS8_2
      port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
            std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal outCarryGen_7_port, outCarryGen_6_port, outCarryGen_5_port, 
      outCarryGen_4_port, outCarryGen_3_port, outCarryGen_2_port, 
      outCarryGen_1_port, outCarryGen_0_port : std_logic;

begin
   
   CG : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Cin => Cin, Co(7) 
                           => outCarryGen_7_port, Co(6) => outCarryGen_6_port, 
                           Co(5) => outCarryGen_5_port, Co(4) => 
                           outCarryGen_4_port, Co(3) => outCarryGen_3_port, 
                           Co(2) => outCarryGen_2_port, Co(1) => 
                           outCarryGen_1_port, Co(0) => outCarryGen_0_port);
   SG : SUMGEN_NBIT32_NBLOCKS8_2 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), cin_vect(7) => 
                           outCarryGen_7_port, cin_vect(6) => 
                           outCarryGen_6_port, cin_vect(5) => 
                           outCarryGen_5_port, cin_vect(4) => 
                           outCarryGen_4_port, cin_vect(3) => 
                           outCarryGen_3_port, cin_vect(2) => 
                           outCarryGen_2_port, cin_vect(1) => 
                           outCarryGen_1_port, cin_vect(0) => 
                           outCarryGen_0_port, Co => Cout, SUM(31) => Y(31), 
                           SUM(30) => Y(30), SUM(29) => Y(29), SUM(28) => Y(28)
                           , SUM(27) => Y(27), SUM(26) => Y(26), SUM(25) => 
                           Y(25), SUM(24) => Y(24), SUM(23) => Y(23), SUM(22) 
                           => Y(22), SUM(21) => Y(21), SUM(20) => Y(20), 
                           SUM(19) => Y(19), SUM(18) => Y(18), SUM(17) => Y(17)
                           , SUM(16) => Y(16), SUM(15) => Y(15), SUM(14) => 
                           Y(14), SUM(13) => Y(13), SUM(12) => Y(12), SUM(11) 
                           => Y(11), SUM(10) => Y(10), SUM(9) => Y(9), SUM(8) 
                           => Y(8), SUM(7) => Y(7), SUM(6) => Y(6), SUM(5) => 
                           Y(5), SUM(4) => Y(4), SUM(3) => Y(3), SUM(2) => Y(2)
                           , SUM(1) => Y(1), SUM(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity P4_ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic;  Y : out std_logic_vector (31 downto 0));

end P4_ADDER_NBIT32_NBIT_PER_BLOCK4_3;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32_NBIT_PER_BLOCK4_3 is

   component SUMGEN_NBIT32_NBLOCKS8_3
      port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
            std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal outCarryGen_7_port, outCarryGen_6_port, outCarryGen_5_port, 
      outCarryGen_4_port, outCarryGen_3_port, outCarryGen_2_port, 
      outCarryGen_1_port, outCarryGen_0_port : std_logic;

begin
   
   CG : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Cin => Cin, Co(7) 
                           => outCarryGen_7_port, Co(6) => outCarryGen_6_port, 
                           Co(5) => outCarryGen_5_port, Co(4) => 
                           outCarryGen_4_port, Co(3) => outCarryGen_3_port, 
                           Co(2) => outCarryGen_2_port, Co(1) => 
                           outCarryGen_1_port, Co(0) => outCarryGen_0_port);
   SG : SUMGEN_NBIT32_NBLOCKS8_3 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), cin_vect(7) => 
                           outCarryGen_7_port, cin_vect(6) => 
                           outCarryGen_6_port, cin_vect(5) => 
                           outCarryGen_5_port, cin_vect(4) => 
                           outCarryGen_4_port, cin_vect(3) => 
                           outCarryGen_3_port, cin_vect(2) => 
                           outCarryGen_2_port, cin_vect(1) => 
                           outCarryGen_1_port, cin_vect(0) => 
                           outCarryGen_0_port, Co => Cout, SUM(31) => Y(31), 
                           SUM(30) => Y(30), SUM(29) => Y(29), SUM(28) => Y(28)
                           , SUM(27) => Y(27), SUM(26) => Y(26), SUM(25) => 
                           Y(25), SUM(24) => Y(24), SUM(23) => Y(23), SUM(22) 
                           => Y(22), SUM(21) => Y(21), SUM(20) => Y(20), 
                           SUM(19) => Y(19), SUM(18) => Y(18), SUM(17) => Y(17)
                           , SUM(16) => Y(16), SUM(15) => Y(15), SUM(14) => 
                           Y(14), SUM(13) => Y(13), SUM(12) => Y(12), SUM(11) 
                           => Y(11), SUM(10) => Y(10), SUM(9) => Y(9), SUM(8) 
                           => Y(8), SUM(7) => Y(7), SUM(6) => Y(6), SUM(5) => 
                           Y(5), SUM(4) => Y(4), SUM(3) => Y(3), SUM(2) => Y(2)
                           , SUM(1) => Y(1), SUM(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_8 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_8;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n52, Q => Q(31), 
                           QN => n148);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n52, Q => Q(30), 
                           QN => n147);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n52, Q => Q(29), 
                           QN => n146);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n52, Q => Q(28), 
                           QN => n145);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n52, Q => Q(27), 
                           QN => n144);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n51, Q => Q(26), 
                           QN => n143);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n51, Q => Q(25),
                           QN => n142);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n51, Q => Q(24),
                           QN => n141);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n51, Q => Q(23),
                           QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n51, Q => Q(22),
                           QN => n139);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n51, Q => Q(21),
                           QN => n138);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n52, Q => Q(20),
                           QN => n137);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n136);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n135);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n52, Q => Q(17),
                           QN => n134);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n133);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n132);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n131);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n50, Q => Q(13),
                           QN => n130);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n50, Q => Q(12),
                           QN => n129);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n50, Q => Q(11),
                           QN => n128);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n50, Q => Q(10),
                           QN => n127);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n50, Q => Q(9), 
                           QN => n126);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n50, Q => Q(8), 
                           QN => n125);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n50, Q => Q(7), 
                           QN => n124);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n50, Q => Q(6), 
                           QN => n123);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n50, Q => Q(5), 
                           QN => n122);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n50, Q => Q(4), 
                           QN => n121);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n50, Q => Q(3), 
                           QN => n120);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n50, Q => Q(2), 
                           QN => n119);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n51, Q => Q(1), 
                           QN => n118);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n52, Q => Q(0), 
                           QN => n117);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n50);
   U5 : BUF_X1 port map( A => RESET_n, Z => n51);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n44);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n146, A2 => n40, B1 => n41, B2 => n55, ZN => 
                           n6);
   U20 : INV_X1 port map( A => D(29), ZN => n55);
   U21 : OAI22_X1 port map( A1 => n117, A2 => n39, B1 => n42, B2 => n116, ZN =>
                           n35);
   U22 : INV_X1 port map( A => D(0), ZN => n116);
   U23 : OAI22_X1 port map( A1 => n118, A2 => n40, B1 => n42, B2 => n115, ZN =>
                           n34);
   U24 : INV_X1 port map( A => D(1), ZN => n115);
   U25 : OAI22_X1 port map( A1 => n143, A2 => n39, B1 => n41, B2 => n58, ZN => 
                           n9);
   U26 : INV_X1 port map( A => D(26), ZN => n58);
   U27 : OAI22_X1 port map( A1 => n144, A2 => n40, B1 => n41, B2 => n57, ZN => 
                           n8);
   U28 : INV_X1 port map( A => D(27), ZN => n57);
   U29 : OAI22_X1 port map( A1 => n145, A2 => n39, B1 => n41, B2 => n56, ZN => 
                           n7);
   U30 : OAI22_X1 port map( A1 => n147, A2 => n40, B1 => n42, B2 => n54, ZN => 
                           n5);
   U31 : INV_X1 port map( A => D(30), ZN => n54);
   U32 : OAI22_X1 port map( A1 => n148, A2 => n39, B1 => n42, B2 => n53, ZN => 
                           n4);
   U33 : INV_X1 port map( A => D(31), ZN => n53);
   U34 : OAI22_X1 port map( A1 => n119, A2 => n40, B1 => n43, B2 => n114, ZN =>
                           n33);
   U35 : INV_X1 port map( A => D(2), ZN => n114);
   U36 : OAI22_X1 port map( A1 => n120, A2 => n40, B1 => n43, B2 => n113, ZN =>
                           n32);
   U37 : INV_X1 port map( A => D(3), ZN => n113);
   U38 : OAI22_X1 port map( A1 => n121, A2 => n40, B1 => n43, B2 => n112, ZN =>
                           n31);
   U39 : INV_X1 port map( A => D(4), ZN => n112);
   U40 : OAI22_X1 port map( A1 => n122, A2 => n40, B1 => n43, B2 => n111, ZN =>
                           n30);
   U41 : INV_X1 port map( A => D(5), ZN => n111);
   U42 : OAI22_X1 port map( A1 => n123, A2 => n40, B1 => n44, B2 => n110, ZN =>
                           n29);
   U43 : INV_X1 port map( A => D(6), ZN => n110);
   U44 : OAI22_X1 port map( A1 => n124, A2 => n40, B1 => n44, B2 => n109, ZN =>
                           n28);
   U45 : INV_X1 port map( A => D(7), ZN => n109);
   U46 : OAI22_X1 port map( A1 => n125, A2 => n40, B1 => n44, B2 => n108, ZN =>
                           n27);
   U47 : INV_X1 port map( A => D(8), ZN => n108);
   U48 : OAI22_X1 port map( A1 => n126, A2 => n40, B1 => n44, B2 => n107, ZN =>
                           n26);
   U49 : INV_X1 port map( A => D(9), ZN => n107);
   U50 : OAI22_X1 port map( A1 => n127, A2 => n40, B1 => n45, B2 => n106, ZN =>
                           n25);
   U51 : INV_X1 port map( A => D(10), ZN => n106);
   U52 : OAI22_X1 port map( A1 => n128, A2 => n40, B1 => n45, B2 => n105, ZN =>
                           n24);
   U53 : INV_X1 port map( A => D(11), ZN => n105);
   U54 : OAI22_X1 port map( A1 => n129, A2 => n40, B1 => n45, B2 => n104, ZN =>
                           n23);
   U55 : INV_X1 port map( A => D(12), ZN => n104);
   U56 : OAI22_X1 port map( A1 => n130, A2 => n40, B1 => n45, B2 => n103, ZN =>
                           n22);
   U57 : INV_X1 port map( A => D(13), ZN => n103);
   U58 : OAI22_X1 port map( A1 => n131, A2 => n39, B1 => n46, B2 => n102, ZN =>
                           n21);
   U59 : INV_X1 port map( A => D(14), ZN => n102);
   U60 : OAI22_X1 port map( A1 => n132, A2 => n39, B1 => n46, B2 => n101, ZN =>
                           n20);
   U61 : INV_X1 port map( A => D(15), ZN => n101);
   U62 : OAI22_X1 port map( A1 => n133, A2 => n39, B1 => n46, B2 => n100, ZN =>
                           n19);
   U63 : INV_X1 port map( A => D(16), ZN => n100);
   U64 : OAI22_X1 port map( A1 => n134, A2 => n39, B1 => n46, B2 => n99, ZN => 
                           n18);
   U65 : INV_X1 port map( A => D(17), ZN => n99);
   U66 : OAI22_X1 port map( A1 => n135, A2 => n39, B1 => n47, B2 => n98, ZN => 
                           n17);
   U67 : INV_X1 port map( A => D(18), ZN => n98);
   U68 : OAI22_X1 port map( A1 => n136, A2 => n39, B1 => n47, B2 => n65, ZN => 
                           n16);
   U69 : OAI22_X1 port map( A1 => n137, A2 => n39, B1 => n47, B2 => n64, ZN => 
                           n15);
   U70 : INV_X1 port map( A => D(20), ZN => n64);
   U71 : OAI22_X1 port map( A1 => n138, A2 => n39, B1 => n47, B2 => n63, ZN => 
                           n14);
   U72 : INV_X1 port map( A => D(21), ZN => n63);
   U73 : OAI22_X1 port map( A1 => n139, A2 => n39, B1 => n48, B2 => n62, ZN => 
                           n13);
   U74 : OAI22_X1 port map( A1 => n140, A2 => n39, B1 => n48, B2 => n61, ZN => 
                           n12);
   U75 : INV_X1 port map( A => D(23), ZN => n61);
   U76 : OAI22_X1 port map( A1 => n141, A2 => n39, B1 => n48, B2 => n60, ZN => 
                           n11);
   U77 : INV_X1 port map( A => D(24), ZN => n60);
   U78 : OAI22_X1 port map( A1 => n142, A2 => n39, B1 => n48, B2 => n59, ZN => 
                           n10);
   U79 : INV_X1 port map( A => D(25), ZN => n59);
   U80 : INV_X1 port map( A => D(28), ZN => n56);
   U81 : INV_X1 port map( A => D(19), ZN => n65);
   U82 : INV_X1 port map( A => D(22), ZN => n62);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_9 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_9;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_9 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, net52311, net52312, net52338, net54370, 
      net54368, net54366, net54364, net54362, net54360, net54356, net54354, 
      net54352, net54350, net54498, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n41, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n43, Q => Q(30), 
                           QN => n67);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n43, Q => Q(29), 
                           QN => n68);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n43, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n43, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n42, Q => Q(26), 
                           QN => n71);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n43, Q => Q(25),
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n42, Q => Q(24),
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n42, Q => Q(23),
                           QN => n74);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n42, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n42, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n43, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n42, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n42, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n43, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n42, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n42, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n42, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n41, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n42, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n41, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n41, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n41, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n41, Q => Q(8), 
                           QN => n89);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n41, Q => Q(7), 
                           QN => n90);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n41, Q => Q(6), 
                           QN => n91);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n41, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n41, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n41, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n41, Q => Q(2), 
                           QN => n95);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n42, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n43, Q => Q(0), 
                           QN => n97);
   U2 : OAI22_X1 port map( A1 => n97, A2 => net54354, B1 => n36, B2 => n37, ZN 
                           => n35);
   U3 : BUF_X1 port map( A => n39, Z => n37);
   U4 : OAI22_X1 port map( A1 => n67, A2 => net54354, B1 => n37, B2 => net52311
                           , ZN => n5);
   U5 : OAI22_X1 port map( A1 => n96, A2 => net54354, B1 => n37, B2 => net52338
                           , ZN => n34);
   U6 : OAI22_X1 port map( A1 => n66, A2 => net54354, B1 => net52312, B2 => n37
                           , ZN => n4);
   U7 : BUF_X1 port map( A => Enable_n, Z => n39);
   U8 : BUF_X1 port map( A => n39, Z => net54356);
   U9 : BUF_X1 port map( A => n39, Z => net54360);
   U10 : INV_X1 port map( A => D(0), ZN => n36);
   U11 : INV_X1 port map( A => n38, ZN => net54354);
   U12 : BUF_X1 port map( A => n40, Z => n38);
   U13 : INV_X1 port map( A => n38, ZN => net54350);
   U14 : INV_X1 port map( A => n38, ZN => net54352);
   U15 : BUF_X1 port map( A => Enable_n, Z => n40);
   U16 : BUF_X1 port map( A => n40, Z => net54368);
   U17 : BUF_X1 port map( A => n40, Z => net54370);
   U18 : BUF_X1 port map( A => Enable_n, Z => net54498);
   U19 : BUF_X1 port map( A => RESET_n, Z => n42);
   U20 : BUF_X1 port map( A => RESET_n, Z => n41);
   U21 : BUF_X1 port map( A => RESET_n, Z => n43);
   U22 : BUF_X1 port map( A => net54498, Z => net54362);
   U23 : BUF_X1 port map( A => net54498, Z => net54366);
   U24 : BUF_X1 port map( A => net54498, Z => net54364);
   U25 : INV_X1 port map( A => D(28), ZN => n103);
   U26 : INV_X1 port map( A => D(30), ZN => net52311);
   U27 : OAI22_X1 port map( A1 => n90, A2 => net54352, B1 => net54362, B2 => 
                           n46, ZN => n28);
   U28 : INV_X1 port map( A => D(7), ZN => n46);
   U29 : OAI22_X1 port map( A1 => n80, A2 => net54350, B1 => net54366, B2 => 
                           n60, ZN => n18);
   U30 : INV_X1 port map( A => D(17), ZN => n60);
   U31 : OAI22_X1 port map( A1 => n95, A2 => net54352, B1 => n45, B2 => 
                           net54360, ZN => n33);
   U32 : INV_X1 port map( A => D(2), ZN => n45);
   U33 : OAI22_X1 port map( A1 => n76, A2 => net54350, B1 => net54368, B2 => 
                           n64, ZN => n14);
   U34 : INV_X1 port map( A => D(21), ZN => n64);
   U35 : OAI22_X1 port map( A1 => n88, A2 => net54352, B1 => net54362, B2 => 
                           n52, ZN => n26);
   U36 : INV_X1 port map( A => D(9), ZN => n52);
   U37 : OAI22_X1 port map( A1 => n83, A2 => net54350, B1 => n55, B2 => 
                           net54366, ZN => n21);
   U38 : INV_X1 port map( A => D(14), ZN => n55);
   U39 : OAI22_X1 port map( A1 => n91, A2 => net54352, B1 => n47, B2 => 
                           net54362, ZN => n29);
   U40 : INV_X1 port map( A => D(6), ZN => n47);
   U41 : OAI22_X1 port map( A1 => n77, A2 => net54350, B1 => net54368, B2 => 
                           n65, ZN => n15);
   U42 : INV_X1 port map( A => D(20), ZN => n65);
   U43 : OAI22_X1 port map( A1 => n93, A2 => net54352, B1 => net54360, B2 => 
                           n49, ZN => n31);
   U44 : INV_X1 port map( A => D(4), ZN => n49);
   U45 : OAI22_X1 port map( A1 => n74, A2 => net54350, B1 => net54370, B2 => 
                           n62, ZN => n12);
   U46 : INV_X1 port map( A => D(23), ZN => n62);
   U47 : OAI22_X1 port map( A1 => n86, A2 => net54352, B1 => net54364, B2 => 
                           n50, ZN => n24);
   U48 : INV_X1 port map( A => D(11), ZN => n50);
   U49 : OAI22_X1 port map( A1 => n79, A2 => net54350, B1 => n59, B2 => 
                           net54368, ZN => n17);
   U50 : INV_X1 port map( A => D(18), ZN => n59);
   U51 : OAI22_X1 port map( A1 => n68, A2 => net54354, B1 => net54356, B2 => 
                           n102, ZN => n6);
   U52 : INV_X1 port map( A => D(29), ZN => n102);
   U53 : INV_X1 port map( A => D(1), ZN => net52338);
   U54 : OAI22_X1 port map( A1 => n82, A2 => net54350, B1 => net54366, B2 => 
                           n54, ZN => n20);
   U55 : INV_X1 port map( A => D(15), ZN => n54);
   U56 : OAI22_X1 port map( A1 => n72, A2 => net54350, B1 => net54370, B2 => 
                           n100, ZN => n10);
   U57 : INV_X1 port map( A => D(25), ZN => n100);
   U58 : OAI22_X1 port map( A1 => n70, A2 => net54354, B1 => net54356, B2 => 
                           n98, ZN => n8);
   U59 : INV_X1 port map( A => D(27), ZN => n98);
   U60 : OAI22_X1 port map( A1 => n71, A2 => net54354, B1 => net54356, B2 => 
                           n99, ZN => n9);
   U61 : INV_X1 port map( A => D(26), ZN => n99);
   U62 : OAI22_X1 port map( A1 => n81, A2 => net54350, B1 => net54366, B2 => 
                           n61, ZN => n19);
   U63 : INV_X1 port map( A => D(16), ZN => n61);
   U64 : OAI22_X1 port map( A1 => n73, A2 => net54350, B1 => net54370, B2 => 
                           n101, ZN => n11);
   U65 : INV_X1 port map( A => D(24), ZN => n101);
   U66 : OAI22_X1 port map( A1 => n87, A2 => net54352, B1 => net54364, B2 => 
                           n51, ZN => n25);
   U67 : INV_X1 port map( A => D(10), ZN => n51);
   U68 : OAI22_X1 port map( A1 => n94, A2 => net54352, B1 => net54360, B2 => 
                           n44, ZN => n32);
   U69 : INV_X1 port map( A => D(3), ZN => n44);
   U70 : OAI22_X1 port map( A1 => n75, A2 => net54350, B1 => net54370, B2 => 
                           n63, ZN => n13);
   U71 : INV_X1 port map( A => D(22), ZN => n63);
   U72 : OAI22_X1 port map( A1 => n78, A2 => net54350, B1 => net54368, B2 => 
                           n58, ZN => n16);
   U73 : INV_X1 port map( A => D(19), ZN => n58);
   U74 : OAI22_X1 port map( A1 => n89, A2 => net54352, B1 => net54362, B2 => 
                           n53, ZN => n27);
   U75 : INV_X1 port map( A => D(8), ZN => n53);
   U76 : OAI22_X1 port map( A1 => n84, A2 => net54352, B1 => net54364, B2 => 
                           n56, ZN => n22);
   U77 : INV_X1 port map( A => D(13), ZN => n56);
   U78 : OAI22_X1 port map( A1 => n69, A2 => net54354, B1 => n103, B2 => 
                           net54356, ZN => n7);
   U79 : INV_X1 port map( A => D(31), ZN => net52312);
   U80 : OAI22_X1 port map( A1 => n85, A2 => net54352, B1 => n57, B2 => 
                           net54364, ZN => n23);
   U81 : INV_X1 port map( A => D(12), ZN => n57);
   U82 : INV_X1 port map( A => D(5), ZN => n48);
   U83 : OAI22_X1 port map( A1 => n92, A2 => net54352, B1 => n48, B2 => 
                           net54360, ZN => n30);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity alu is

   port( data_in1, data_in2 : in std_logic_vector (31 downto 0);  op_sel : in 
         std_logic_vector (3 downto 0);  data_out : out std_logic_vector (31 
         downto 0));

end alu;

architecture SYN_BEH of alu is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component mux11to1_nbit32
      port( A, B, C, D, E, F, H : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (3 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component comparator
      port( r1, r2 : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (2 downto 0);  data_out : out std_logic_vector (31
            downto 0));
   end component;
   
   component shifter_dx_nbit32
      port( r1, r2 : in std_logic_vector (31 downto 0);  log : in std_logic;  
            data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component shifter_sx_nbit32
      port( r1, r2 : in std_logic_vector (31 downto 0);  data_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component xor_gate_nbit32
      port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component or_gate_nbit32
      port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component and_gate_nbit32
      port( A, B : in std_logic_vector (31 downto 0);  Y : out std_logic_vector
            (31 downto 0));
   end component;
   
   component P4_ADDER_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal p4_cin, add_sel, mux_sel_3_port, mux_sel_2_port, mux_sel_1_port, 
      mux_sel_0_port, log_shift, cmp_sel_2_port, cmp_sel_1_port, cmp_sel_0_port
      , N41, N42, N43, N44, N49, p4_operand_31_port, p4_operand_30_port, 
      p4_operand_29_port, p4_operand_28_port, p4_operand_27_port, 
      p4_operand_26_port, p4_operand_25_port, p4_operand_24_port, 
      p4_operand_23_port, p4_operand_22_port, p4_operand_21_port, 
      p4_operand_20_port, p4_operand_19_port, p4_operand_18_port, 
      p4_operand_17_port, p4_operand_16_port, p4_operand_15_port, 
      p4_operand_14_port, p4_operand_13_port, p4_operand_12_port, 
      p4_operand_11_port, p4_operand_10_port, p4_operand_9_port, 
      p4_operand_8_port, p4_operand_7_port, p4_operand_6_port, 
      p4_operand_5_port, p4_operand_4_port, p4_operand_3_port, 
      p4_operand_2_port, p4_operand_1_port, p4_operand_0_port, p4_out_31_port, 
      p4_out_30_port, p4_out_29_port, p4_out_28_port, p4_out_27_port, 
      p4_out_26_port, p4_out_25_port, p4_out_24_port, p4_out_23_port, 
      p4_out_22_port, p4_out_21_port, p4_out_20_port, p4_out_19_port, 
      p4_out_18_port, p4_out_17_port, p4_out_16_port, p4_out_15_port, 
      p4_out_14_port, p4_out_13_port, p4_out_12_port, p4_out_11_port, 
      p4_out_10_port, p4_out_9_port, p4_out_8_port, p4_out_7_port, 
      p4_out_6_port, p4_out_5_port, p4_out_4_port, p4_out_3_port, p4_out_2_port
      , p4_out_1_port, p4_out_0_port, and_out_31_port, and_out_30_port, 
      and_out_29_port, and_out_28_port, and_out_27_port, and_out_26_port, 
      and_out_25_port, and_out_24_port, and_out_23_port, and_out_22_port, 
      and_out_21_port, and_out_20_port, and_out_19_port, and_out_18_port, 
      and_out_17_port, and_out_16_port, and_out_15_port, and_out_14_port, 
      and_out_13_port, and_out_12_port, and_out_11_port, and_out_10_port, 
      and_out_9_port, and_out_8_port, and_out_7_port, and_out_6_port, 
      and_out_5_port, and_out_4_port, and_out_3_port, and_out_2_port, 
      and_out_1_port, and_out_0_port, or_out_31_port, or_out_30_port, 
      or_out_29_port, or_out_28_port, or_out_27_port, or_out_26_port, 
      or_out_25_port, or_out_24_port, or_out_23_port, or_out_22_port, 
      or_out_21_port, or_out_20_port, or_out_19_port, or_out_18_port, 
      or_out_17_port, or_out_16_port, or_out_15_port, or_out_14_port, 
      or_out_13_port, or_out_12_port, or_out_11_port, or_out_10_port, 
      or_out_9_port, or_out_8_port, or_out_7_port, or_out_6_port, or_out_5_port
      , or_out_4_port, or_out_3_port, or_out_2_port, or_out_1_port, 
      or_out_0_port, xor_out_31_port, xor_out_30_port, xor_out_29_port, 
      xor_out_28_port, xor_out_27_port, xor_out_26_port, xor_out_25_port, 
      xor_out_24_port, xor_out_23_port, xor_out_22_port, xor_out_21_port, 
      xor_out_20_port, xor_out_19_port, xor_out_18_port, xor_out_17_port, 
      xor_out_16_port, xor_out_15_port, xor_out_14_port, xor_out_13_port, 
      xor_out_12_port, xor_out_11_port, xor_out_10_port, xor_out_9_port, 
      xor_out_8_port, xor_out_7_port, xor_out_6_port, xor_out_5_port, 
      xor_out_4_port, xor_out_3_port, xor_out_2_port, xor_out_1_port, 
      xor_out_0_port, sl_out_31_port, sl_out_30_port, sl_out_29_port, 
      sl_out_28_port, sl_out_27_port, sl_out_26_port, sl_out_25_port, 
      sl_out_24_port, sl_out_23_port, sl_out_22_port, sl_out_21_port, 
      sl_out_20_port, sl_out_19_port, sl_out_18_port, sl_out_17_port, 
      sl_out_16_port, sl_out_15_port, sl_out_14_port, sl_out_13_port, 
      sl_out_12_port, sl_out_11_port, sl_out_10_port, sl_out_9_port, 
      sl_out_8_port, sl_out_7_port, sl_out_6_port, sl_out_5_port, sl_out_4_port
      , sl_out_3_port, sl_out_2_port, sl_out_1_port, sl_out_0_port, 
      sr_out_31_port, sr_out_30_port, sr_out_29_port, sr_out_28_port, 
      sr_out_27_port, sr_out_26_port, sr_out_25_port, sr_out_24_port, 
      sr_out_23_port, sr_out_22_port, sr_out_21_port, sr_out_20_port, 
      sr_out_19_port, sr_out_18_port, sr_out_17_port, sr_out_16_port, 
      sr_out_15_port, sr_out_14_port, sr_out_13_port, sr_out_12_port, 
      sr_out_11_port, sr_out_10_port, sr_out_9_port, sr_out_8_port, 
      sr_out_7_port, sr_out_6_port, sr_out_5_port, sr_out_4_port, sr_out_3_port
      , sr_out_2_port, sr_out_1_port, sr_out_0_port, cmp_out_31_port, 
      cmp_out_30_port, cmp_out_29_port, cmp_out_28_port, cmp_out_27_port, 
      cmp_out_26_port, cmp_out_25_port, cmp_out_24_port, cmp_out_23_port, 
      cmp_out_22_port, cmp_out_21_port, cmp_out_20_port, cmp_out_19_port, 
      cmp_out_18_port, cmp_out_17_port, cmp_out_16_port, cmp_out_15_port, 
      cmp_out_14_port, cmp_out_13_port, cmp_out_12_port, cmp_out_11_port, 
      cmp_out_10_port, cmp_out_9_port, cmp_out_8_port, cmp_out_7_port, 
      cmp_out_6_port, cmp_out_5_port, cmp_out_4_port, cmp_out_3_port, 
      cmp_out_2_port, cmp_out_1_port, cmp_out_0_port, n54, n55, n56, n40, 
      n41_port, n42_port, n43_port, n44_port, n45, n46, n47, n48, n49_port, n50
      , n51, n52, n53, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197 : std_logic;

begin
   
   cmp_sel_reg_2_inst : DLH_X1 port map( G => n121, D => N49, Q => 
                           cmp_sel_2_port);
   cmp_sel_reg_1_inst : DLH_X1 port map( G => n121, D => n55, Q => 
                           cmp_sel_1_port);
   cmp_sel_reg_0_inst : DLH_X1 port map( G => n121, D => n54, Q => 
                           cmp_sel_0_port);
   p4_cin_reg : DLH_X1 port map( G => N41, D => n56, Q => p4_cin);
   mux_sel_reg_2_inst : DLH_X1 port map( G => N42, D => n50, Q => 
                           mux_sel_2_port);
   mux_sel_reg_1_inst : DLH_X1 port map( G => N42, D => N44, Q => 
                           mux_sel_1_port);
   mux_sel_reg_0_inst : DLH_X1 port map( G => N42, D => N43, Q => 
                           mux_sel_0_port);
   log_shift_reg : DLH_X1 port map( G => n123, D => n51, Q => log_shift);
   mux_sel_3_port <= '0';
   cmp_out_1_port <= '0';
   cmp_out_2_port <= '0';
   cmp_out_3_port <= '0';
   cmp_out_4_port <= '0';
   cmp_out_5_port <= '0';
   cmp_out_6_port <= '0';
   cmp_out_7_port <= '0';
   cmp_out_8_port <= '0';
   cmp_out_9_port <= '0';
   cmp_out_10_port <= '0';
   cmp_out_11_port <= '0';
   cmp_out_12_port <= '0';
   cmp_out_13_port <= '0';
   cmp_out_14_port <= '0';
   cmp_out_15_port <= '0';
   cmp_out_16_port <= '0';
   cmp_out_17_port <= '0';
   cmp_out_18_port <= '0';
   cmp_out_19_port <= '0';
   cmp_out_20_port <= '0';
   cmp_out_21_port <= '0';
   cmp_out_22_port <= '0';
   cmp_out_23_port <= '0';
   cmp_out_24_port <= '0';
   cmp_out_25_port <= '0';
   cmp_out_26_port <= '0';
   cmp_out_27_port <= '0';
   cmp_out_28_port <= '0';
   cmp_out_29_port <= '0';
   cmp_out_30_port <= '0';
   cmp_out_31_port <= '0';
   U57 : NAND3_X1 port map( A1 => n42_port, A2 => n40, A3 => n43_port, ZN => 
                           N44);
   U58 : NAND3_X1 port map( A1 => n42_port, A2 => n122, A3 => n44_port, ZN => 
                           N42);
   U59 : XOR2_X1 port map( A => op_sel(2), B => op_sel(0), Z => n46);
   U60 : XOR2_X1 port map( A => op_sel(1), B => op_sel(0), Z => n49_port);
   U61 : NAND3_X1 port map( A1 => n127, A2 => n126, A3 => op_sel(2), ZN => 
                           n42_port);
   mux_p4 : MUX21_GENERIC_NBIT32_2 port map( A(31) => data_in2(31), A(30) => 
                           n61, A(29) => n78, A(28) => n64, A(27) => 
                           data_in2(27), A(26) => n62, A(25) => data_in2(25), 
                           A(24) => n52, A(23) => n60, A(22) => n57, A(21) => 
                           n75, A(20) => data_in2(20), A(19) => n73, A(18) => 
                           data_in2(18), A(17) => data_in2(17), A(16) => 
                           data_in2(16), A(15) => data_in2(15), A(14) => 
                           data_in2(14), A(13) => n53, A(12) => data_in2(12), 
                           A(11) => data_in2(11), A(10) => n58, A(9) => n77, 
                           A(8) => n76, A(7) => n59, A(6) => n74, A(5) => 
                           data_in2(5), A(4) => data_in2(4), A(3) => n63, A(2) 
                           => n70, A(1) => n68, A(0) => n72, B(31) => n89, 
                           B(30) => n90, B(29) => n91, B(28) => n92, B(27) => 
                           n93, B(26) => n94, B(25) => n95, B(24) => n96, B(23)
                           => n97, B(22) => n98, B(21) => n99, B(20) => n100, 
                           B(19) => n101, B(18) => n102, B(17) => n103, B(16) 
                           => n104, B(15) => n105, B(14) => n106, B(13) => n107
                           , B(12) => n108, B(11) => n109, B(10) => n110, B(9) 
                           => n111, B(8) => n112, B(7) => n113, B(6) => n114, 
                           B(5) => n115, B(4) => n116, B(3) => n117, B(2) => 
                           n118, B(1) => n119, B(0) => n120, SEL => add_sel, 
                           Y(31) => p4_operand_31_port, Y(30) => 
                           p4_operand_30_port, Y(29) => p4_operand_29_port, 
                           Y(28) => p4_operand_28_port, Y(27) => 
                           p4_operand_27_port, Y(26) => p4_operand_26_port, 
                           Y(25) => p4_operand_25_port, Y(24) => 
                           p4_operand_24_port, Y(23) => p4_operand_23_port, 
                           Y(22) => p4_operand_22_port, Y(21) => 
                           p4_operand_21_port, Y(20) => p4_operand_20_port, 
                           Y(19) => p4_operand_19_port, Y(18) => 
                           p4_operand_18_port, Y(17) => p4_operand_17_port, 
                           Y(16) => p4_operand_16_port, Y(15) => 
                           p4_operand_15_port, Y(14) => p4_operand_14_port, 
                           Y(13) => p4_operand_13_port, Y(12) => 
                           p4_operand_12_port, Y(11) => p4_operand_11_port, 
                           Y(10) => p4_operand_10_port, Y(9) => 
                           p4_operand_9_port, Y(8) => p4_operand_8_port, Y(7) 
                           => p4_operand_7_port, Y(6) => p4_operand_6_port, 
                           Y(5) => p4_operand_5_port, Y(4) => p4_operand_4_port
                           , Y(3) => p4_operand_3_port, Y(2) => 
                           p4_operand_2_port, Y(1) => p4_operand_1_port, Y(0) 
                           => p4_operand_0_port);
   add : P4_ADDER_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => data_in1(31), 
                           A(30) => n88, A(29) => data_in1(29), A(28) => 
                           data_in1(28), A(27) => data_in1(27), A(26) => 
                           data_in1(26), A(25) => data_in1(25), A(24) => 
                           data_in1(24), A(23) => data_in1(23), A(22) => n87, 
                           A(21) => n86, A(20) => data_in1(20), A(19) => 
                           data_in1(19), A(18) => n85, A(17) => data_in1(17), 
                           A(16) => data_in1(16), A(15) => data_in1(15), A(14) 
                           => n84, A(13) => n83, A(12) => data_in1(12), A(11) 
                           => data_in1(11), A(10) => data_in1(10), A(9) => n82,
                           A(8) => n81, A(7) => data_in1(7), A(6) => 
                           data_in1(6), A(5) => data_in1(5), A(4) => n80, A(3) 
                           => data_in1(3), A(2) => n67, A(1) => n66, A(0) => 
                           n79, B(31) => p4_operand_31_port, B(30) => 
                           p4_operand_30_port, B(29) => p4_operand_29_port, 
                           B(28) => p4_operand_28_port, B(27) => 
                           p4_operand_27_port, B(26) => p4_operand_26_port, 
                           B(25) => p4_operand_25_port, B(24) => 
                           p4_operand_24_port, B(23) => p4_operand_23_port, 
                           B(22) => p4_operand_22_port, B(21) => 
                           p4_operand_21_port, B(20) => p4_operand_20_port, 
                           B(19) => p4_operand_19_port, B(18) => 
                           p4_operand_18_port, B(17) => p4_operand_17_port, 
                           B(16) => p4_operand_16_port, B(15) => 
                           p4_operand_15_port, B(14) => p4_operand_14_port, 
                           B(13) => p4_operand_13_port, B(12) => 
                           p4_operand_12_port, B(11) => p4_operand_11_port, 
                           B(10) => p4_operand_10_port, B(9) => 
                           p4_operand_9_port, B(8) => p4_operand_8_port, B(7) 
                           => p4_operand_7_port, B(6) => p4_operand_6_port, 
                           B(5) => p4_operand_5_port, B(4) => p4_operand_4_port
                           , B(3) => p4_operand_3_port, B(2) => 
                           p4_operand_2_port, B(1) => p4_operand_1_port, B(0) 
                           => p4_operand_0_port, Cin => p4_cin, Cout => n_1166,
                           Y(31) => p4_out_31_port, Y(30) => p4_out_30_port, 
                           Y(29) => p4_out_29_port, Y(28) => p4_out_28_port, 
                           Y(27) => p4_out_27_port, Y(26) => p4_out_26_port, 
                           Y(25) => p4_out_25_port, Y(24) => p4_out_24_port, 
                           Y(23) => p4_out_23_port, Y(22) => p4_out_22_port, 
                           Y(21) => p4_out_21_port, Y(20) => p4_out_20_port, 
                           Y(19) => p4_out_19_port, Y(18) => p4_out_18_port, 
                           Y(17) => p4_out_17_port, Y(16) => p4_out_16_port, 
                           Y(15) => p4_out_15_port, Y(14) => p4_out_14_port, 
                           Y(13) => p4_out_13_port, Y(12) => p4_out_12_port, 
                           Y(11) => p4_out_11_port, Y(10) => p4_out_10_port, 
                           Y(9) => p4_out_9_port, Y(8) => p4_out_8_port, Y(7) 
                           => p4_out_7_port, Y(6) => p4_out_6_port, Y(5) => 
                           p4_out_5_port, Y(4) => p4_out_4_port, Y(3) => 
                           p4_out_3_port, Y(2) => p4_out_2_port, Y(1) => 
                           p4_out_1_port, Y(0) => p4_out_0_port);
   and_m : and_gate_nbit32 port map( A(31) => data_in1(31), A(30) => n88, A(29)
                           => data_in1(29), A(28) => data_in1(28), A(27) => 
                           data_in1(27), A(26) => data_in1(26), A(25) => 
                           data_in1(25), A(24) => data_in1(24), A(23) => 
                           data_in1(23), A(22) => n87, A(21) => n86, A(20) => 
                           data_in1(20), A(19) => data_in1(19), A(18) => n85, 
                           A(17) => data_in1(17), A(16) => data_in1(16), A(15) 
                           => data_in1(15), A(14) => n84, A(13) => n83, A(12) 
                           => data_in1(12), A(11) => data_in1(11), A(10) => 
                           data_in1(10), A(9) => n82, A(8) => n81, A(7) => 
                           data_in1(7), A(6) => data_in1(6), A(5) => 
                           data_in1(5), A(4) => n80, A(3) => data_in1(3), A(2) 
                           => n67, A(1) => n66, A(0) => n79, B(31) => 
                           data_in2(31), B(30) => n61, B(29) => n78, B(28) => 
                           n64, B(27) => data_in2(27), B(26) => n62, B(25) => 
                           data_in2(25), B(24) => n52, B(23) => n60, B(22) => 
                           n57, B(21) => n75, B(20) => data_in2(20), B(19) => 
                           n73, B(18) => data_in2(18), B(17) => data_in2(17), 
                           B(16) => data_in2(16), B(15) => data_in2(15), B(14) 
                           => data_in2(14), B(13) => n53, B(12) => data_in2(12)
                           , B(11) => data_in2(11), B(10) => n58, B(9) => n77, 
                           B(8) => n76, B(7) => n59, B(6) => n74, B(5) => 
                           data_in2(5), B(4) => data_in2(4), B(3) => n63, B(2) 
                           => n71, B(1) => n69, B(0) => n72, Y(31) => 
                           and_out_31_port, Y(30) => and_out_30_port, Y(29) => 
                           and_out_29_port, Y(28) => and_out_28_port, Y(27) => 
                           and_out_27_port, Y(26) => and_out_26_port, Y(25) => 
                           and_out_25_port, Y(24) => and_out_24_port, Y(23) => 
                           and_out_23_port, Y(22) => and_out_22_port, Y(21) => 
                           and_out_21_port, Y(20) => and_out_20_port, Y(19) => 
                           and_out_19_port, Y(18) => and_out_18_port, Y(17) => 
                           and_out_17_port, Y(16) => and_out_16_port, Y(15) => 
                           and_out_15_port, Y(14) => and_out_14_port, Y(13) => 
                           and_out_13_port, Y(12) => and_out_12_port, Y(11) => 
                           and_out_11_port, Y(10) => and_out_10_port, Y(9) => 
                           and_out_9_port, Y(8) => and_out_8_port, Y(7) => 
                           and_out_7_port, Y(6) => and_out_6_port, Y(5) => 
                           and_out_5_port, Y(4) => and_out_4_port, Y(3) => 
                           and_out_3_port, Y(2) => and_out_2_port, Y(1) => 
                           and_out_1_port, Y(0) => and_out_0_port);
   or_m : or_gate_nbit32 port map( A(31) => data_in1(31), A(30) => n88, A(29) 
                           => data_in1(29), A(28) => data_in1(28), A(27) => 
                           data_in1(27), A(26) => data_in1(26), A(25) => 
                           data_in1(25), A(24) => data_in1(24), A(23) => 
                           data_in1(23), A(22) => n87, A(21) => n86, A(20) => 
                           data_in1(20), A(19) => data_in1(19), A(18) => n85, 
                           A(17) => data_in1(17), A(16) => data_in1(16), A(15) 
                           => data_in1(15), A(14) => n84, A(13) => n83, A(12) 
                           => data_in1(12), A(11) => data_in1(11), A(10) => 
                           data_in1(10), A(9) => n82, A(8) => n81, A(7) => 
                           data_in1(7), A(6) => data_in1(6), A(5) => 
                           data_in1(5), A(4) => n80, A(3) => data_in1(3), A(2) 
                           => n67, A(1) => n66, A(0) => n79, B(31) => 
                           data_in2(31), B(30) => n61, B(29) => n78, B(28) => 
                           n64, B(27) => data_in2(27), B(26) => n62, B(25) => 
                           data_in2(25), B(24) => n52, B(23) => n60, B(22) => 
                           n57, B(21) => n75, B(20) => data_in2(20), B(19) => 
                           n73, B(18) => data_in2(18), B(17) => data_in2(17), 
                           B(16) => data_in2(16), B(15) => data_in2(15), B(14) 
                           => data_in2(14), B(13) => n53, B(12) => data_in2(12)
                           , B(11) => data_in2(11), B(10) => n58, B(9) => n77, 
                           B(8) => n76, B(7) => n59, B(6) => n74, B(5) => 
                           data_in2(5), B(4) => data_in2(4), B(3) => n63, B(2) 
                           => n71, B(1) => n69, B(0) => n72, Y(31) => 
                           or_out_31_port, Y(30) => or_out_30_port, Y(29) => 
                           or_out_29_port, Y(28) => or_out_28_port, Y(27) => 
                           or_out_27_port, Y(26) => or_out_26_port, Y(25) => 
                           or_out_25_port, Y(24) => or_out_24_port, Y(23) => 
                           or_out_23_port, Y(22) => or_out_22_port, Y(21) => 
                           or_out_21_port, Y(20) => or_out_20_port, Y(19) => 
                           or_out_19_port, Y(18) => or_out_18_port, Y(17) => 
                           or_out_17_port, Y(16) => or_out_16_port, Y(15) => 
                           or_out_15_port, Y(14) => or_out_14_port, Y(13) => 
                           or_out_13_port, Y(12) => or_out_12_port, Y(11) => 
                           or_out_11_port, Y(10) => or_out_10_port, Y(9) => 
                           or_out_9_port, Y(8) => or_out_8_port, Y(7) => 
                           or_out_7_port, Y(6) => or_out_6_port, Y(5) => 
                           or_out_5_port, Y(4) => or_out_4_port, Y(3) => 
                           or_out_3_port, Y(2) => or_out_2_port, Y(1) => 
                           or_out_1_port, Y(0) => or_out_0_port);
   xor_m : xor_gate_nbit32 port map( A(31) => data_in1(31), A(30) => n88, A(29)
                           => data_in1(29), A(28) => data_in1(28), A(27) => 
                           data_in1(27), A(26) => data_in1(26), A(25) => 
                           data_in1(25), A(24) => data_in1(24), A(23) => 
                           data_in1(23), A(22) => n87, A(21) => n86, A(20) => 
                           data_in1(20), A(19) => data_in1(19), A(18) => n85, 
                           A(17) => data_in1(17), A(16) => data_in1(16), A(15) 
                           => data_in1(15), A(14) => n84, A(13) => n83, A(12) 
                           => data_in1(12), A(11) => data_in1(11), A(10) => 
                           data_in1(10), A(9) => n82, A(8) => n81, A(7) => 
                           data_in1(7), A(6) => data_in1(6), A(5) => 
                           data_in1(5), A(4) => n80, A(3) => data_in1(3), A(2) 
                           => n67, A(1) => n66, A(0) => n79, B(31) => 
                           data_in2(31), B(30) => n61, B(29) => n78, B(28) => 
                           n64, B(27) => data_in2(27), B(26) => n62, B(25) => 
                           data_in2(25), B(24) => n52, B(23) => n60, B(22) => 
                           n57, B(21) => n75, B(20) => data_in2(20), B(19) => 
                           n73, B(18) => data_in2(18), B(17) => data_in2(17), 
                           B(16) => data_in2(16), B(15) => data_in2(15), B(14) 
                           => data_in2(14), B(13) => n53, B(12) => data_in2(12)
                           , B(11) => data_in2(11), B(10) => n58, B(9) => n77, 
                           B(8) => n76, B(7) => n59, B(6) => n74, B(5) => 
                           data_in2(5), B(4) => data_in2(4), B(3) => n63, B(2) 
                           => n70, B(1) => n68, B(0) => n72, Y(31) => 
                           xor_out_31_port, Y(30) => xor_out_30_port, Y(29) => 
                           xor_out_29_port, Y(28) => xor_out_28_port, Y(27) => 
                           xor_out_27_port, Y(26) => xor_out_26_port, Y(25) => 
                           xor_out_25_port, Y(24) => xor_out_24_port, Y(23) => 
                           xor_out_23_port, Y(22) => xor_out_22_port, Y(21) => 
                           xor_out_21_port, Y(20) => xor_out_20_port, Y(19) => 
                           xor_out_19_port, Y(18) => xor_out_18_port, Y(17) => 
                           xor_out_17_port, Y(16) => xor_out_16_port, Y(15) => 
                           xor_out_15_port, Y(14) => xor_out_14_port, Y(13) => 
                           xor_out_13_port, Y(12) => xor_out_12_port, Y(11) => 
                           xor_out_11_port, Y(10) => xor_out_10_port, Y(9) => 
                           xor_out_9_port, Y(8) => xor_out_8_port, Y(7) => 
                           xor_out_7_port, Y(6) => xor_out_6_port, Y(5) => 
                           xor_out_5_port, Y(4) => xor_out_4_port, Y(3) => 
                           xor_out_3_port, Y(2) => xor_out_2_port, Y(1) => 
                           xor_out_1_port, Y(0) => xor_out_0_port);
   sl : shifter_sx_nbit32 port map( r1(31) => data_in1(31), r1(30) => n88, 
                           r1(29) => data_in1(29), r1(28) => data_in1(28), 
                           r1(27) => data_in1(27), r1(26) => data_in1(26), 
                           r1(25) => data_in1(25), r1(24) => data_in1(24), 
                           r1(23) => data_in1(23), r1(22) => n87, r1(21) => n86
                           , r1(20) => data_in1(20), r1(19) => data_in1(19), 
                           r1(18) => n85, r1(17) => data_in1(17), r1(16) => 
                           data_in1(16), r1(15) => data_in1(15), r1(14) => n84,
                           r1(13) => n83, r1(12) => data_in1(12), r1(11) => 
                           data_in1(11), r1(10) => data_in1(10), r1(9) => n82, 
                           r1(8) => n81, r1(7) => data_in1(7), r1(6) => 
                           data_in1(6), r1(5) => data_in1(5), r1(4) => n80, 
                           r1(3) => data_in1(3), r1(2) => n67, r1(1) => n66, 
                           r1(0) => n79, r2(31) => data_in2(31), r2(30) => 
                           data_in2(30), r2(29) => data_in2(29), r2(28) => 
                           data_in2(28), r2(27) => data_in2(27), r2(26) => 
                           data_in2(26), r2(25) => data_in2(25), r2(24) => 
                           data_in2(24), r2(23) => data_in2(23), r2(22) => 
                           data_in2(22), r2(21) => data_in2(21), r2(20) => 
                           data_in2(20), r2(19) => data_in2(19), r2(18) => 
                           data_in2(18), r2(17) => data_in2(17), r2(16) => 
                           data_in2(16), r2(15) => data_in2(15), r2(14) => 
                           data_in2(14), r2(13) => data_in2(13), r2(12) => 
                           data_in2(12), r2(11) => data_in2(11), r2(10) => 
                           data_in2(10), r2(9) => data_in2(9), r2(8) => 
                           data_in2(8), r2(7) => data_in2(7), r2(6) => 
                           data_in2(6), r2(5) => data_in2(5), r2(4) => 
                           data_in2(4), r2(3) => n63, r2(2) => n71, r2(1) => 
                           n69, r2(0) => n72, data_out(31) => sl_out_31_port, 
                           data_out(30) => sl_out_30_port, data_out(29) => 
                           sl_out_29_port, data_out(28) => sl_out_28_port, 
                           data_out(27) => sl_out_27_port, data_out(26) => 
                           sl_out_26_port, data_out(25) => sl_out_25_port, 
                           data_out(24) => sl_out_24_port, data_out(23) => 
                           sl_out_23_port, data_out(22) => sl_out_22_port, 
                           data_out(21) => sl_out_21_port, data_out(20) => 
                           sl_out_20_port, data_out(19) => sl_out_19_port, 
                           data_out(18) => sl_out_18_port, data_out(17) => 
                           sl_out_17_port, data_out(16) => sl_out_16_port, 
                           data_out(15) => sl_out_15_port, data_out(14) => 
                           sl_out_14_port, data_out(13) => sl_out_13_port, 
                           data_out(12) => sl_out_12_port, data_out(11) => 
                           sl_out_11_port, data_out(10) => sl_out_10_port, 
                           data_out(9) => sl_out_9_port, data_out(8) => 
                           sl_out_8_port, data_out(7) => sl_out_7_port, 
                           data_out(6) => sl_out_6_port, data_out(5) => 
                           sl_out_5_port, data_out(4) => sl_out_4_port, 
                           data_out(3) => sl_out_3_port, data_out(2) => 
                           sl_out_2_port, data_out(1) => sl_out_1_port, 
                           data_out(0) => sl_out_0_port);
   sr : shifter_dx_nbit32 port map( r1(31) => data_in1(31), r1(30) => n88, 
                           r1(29) => data_in1(29), r1(28) => data_in1(28), 
                           r1(27) => data_in1(27), r1(26) => data_in1(26), 
                           r1(25) => data_in1(25), r1(24) => data_in1(24), 
                           r1(23) => data_in1(23), r1(22) => n87, r1(21) => n86
                           , r1(20) => data_in1(20), r1(19) => data_in1(19), 
                           r1(18) => n85, r1(17) => data_in1(17), r1(16) => 
                           data_in1(16), r1(15) => data_in1(15), r1(14) => n84,
                           r1(13) => n83, r1(12) => data_in1(12), r1(11) => 
                           data_in1(11), r1(10) => data_in1(10), r1(9) => n82, 
                           r1(8) => n81, r1(7) => data_in1(7), r1(6) => 
                           data_in1(6), r1(5) => data_in1(5), r1(4) => n80, 
                           r1(3) => data_in1(3), r1(2) => n67, r1(1) => n66, 
                           r1(0) => n79, r2(31) => data_in2(31), r2(30) => n61,
                           r2(29) => data_in2(29), r2(28) => data_in2(28), 
                           r2(27) => data_in2(27), r2(26) => data_in2(26), 
                           r2(25) => data_in2(25), r2(24) => data_in2(24), 
                           r2(23) => data_in2(23), r2(22) => data_in2(22), 
                           r2(21) => data_in2(21), r2(20) => data_in2(20), 
                           r2(19) => data_in2(19), r2(18) => data_in2(18), 
                           r2(17) => data_in2(17), r2(16) => data_in2(16), 
                           r2(15) => data_in2(15), r2(14) => data_in2(14), 
                           r2(13) => data_in2(13), r2(12) => data_in2(12), 
                           r2(11) => data_in2(11), r2(10) => n58, r2(9) => 
                           data_in2(9), r2(8) => data_in2(8), r2(7) => 
                           data_in2(7), r2(6) => data_in2(6), r2(5) => 
                           data_in2(5), r2(4) => data_in2(4), r2(3) => n63, 
                           r2(2) => n70, r2(1) => n68, r2(0) => n72, log => 
                           log_shift, data_out(31) => sr_out_31_port, 
                           data_out(30) => sr_out_30_port, data_out(29) => 
                           sr_out_29_port, data_out(28) => sr_out_28_port, 
                           data_out(27) => sr_out_27_port, data_out(26) => 
                           sr_out_26_port, data_out(25) => sr_out_25_port, 
                           data_out(24) => sr_out_24_port, data_out(23) => 
                           sr_out_23_port, data_out(22) => sr_out_22_port, 
                           data_out(21) => sr_out_21_port, data_out(20) => 
                           sr_out_20_port, data_out(19) => sr_out_19_port, 
                           data_out(18) => sr_out_18_port, data_out(17) => 
                           sr_out_17_port, data_out(16) => sr_out_16_port, 
                           data_out(15) => sr_out_15_port, data_out(14) => 
                           sr_out_14_port, data_out(13) => sr_out_13_port, 
                           data_out(12) => sr_out_12_port, data_out(11) => 
                           sr_out_11_port, data_out(10) => sr_out_10_port, 
                           data_out(9) => sr_out_9_port, data_out(8) => 
                           sr_out_8_port, data_out(7) => sr_out_7_port, 
                           data_out(6) => sr_out_6_port, data_out(5) => 
                           sr_out_5_port, data_out(4) => sr_out_4_port, 
                           data_out(3) => sr_out_3_port, data_out(2) => 
                           sr_out_2_port, data_out(1) => sr_out_1_port, 
                           data_out(0) => sr_out_0_port);
   cmp : comparator port map( r1(31) => data_in1(31), r1(30) => n88, r1(29) => 
                           data_in1(29), r1(28) => data_in1(28), r1(27) => 
                           data_in1(27), r1(26) => data_in1(26), r1(25) => 
                           data_in1(25), r1(24) => data_in1(24), r1(23) => 
                           data_in1(23), r1(22) => n87, r1(21) => n86, r1(20) 
                           => data_in1(20), r1(19) => data_in1(19), r1(18) => 
                           n85, r1(17) => data_in1(17), r1(16) => data_in1(16),
                           r1(15) => data_in1(15), r1(14) => n84, r1(13) => n83
                           , r1(12) => data_in1(12), r1(11) => data_in1(11), 
                           r1(10) => data_in1(10), r1(9) => n82, r1(8) => n81, 
                           r1(7) => data_in1(7), r1(6) => data_in1(6), r1(5) =>
                           data_in1(5), r1(4) => n80, r1(3) => data_in1(3), 
                           r1(2) => data_in1(2), r1(1) => data_in1(1), r1(0) =>
                           data_in1(0), r2(31) => data_in2(31), r2(30) => n61, 
                           r2(29) => n78, r2(28) => n64, r2(27) => data_in2(27)
                           , r2(26) => n62, r2(25) => data_in2(25), r2(24) => 
                           n52, r2(23) => n60, r2(22) => n57, r2(21) => n75, 
                           r2(20) => data_in2(20), r2(19) => n73, r2(18) => 
                           data_in2(18), r2(17) => data_in2(17), r2(16) => 
                           data_in2(16), r2(15) => data_in2(15), r2(14) => 
                           data_in2(14), r2(13) => n53, r2(12) => data_in2(12),
                           r2(11) => data_in2(11), r2(10) => n58, r2(9) => n77,
                           r2(8) => n76, r2(7) => n59, r2(6) => n74, r2(5) => 
                           data_in2(5), r2(4) => data_in2(4), r2(3) => 
                           data_in2(3), r2(2) => data_in2(2), r2(1) => 
                           data_in2(1), r2(0) => data_in2(0), sel(2) => 
                           cmp_sel_2_port, sel(1) => cmp_sel_1_port, sel(0) => 
                           cmp_sel_0_port, data_out(31) => n_1167, data_out(30)
                           => n_1168, data_out(29) => n_1169, data_out(28) => 
                           n_1170, data_out(27) => n_1171, data_out(26) => 
                           n_1172, data_out(25) => n_1173, data_out(24) => 
                           n_1174, data_out(23) => n_1175, data_out(22) => 
                           n_1176, data_out(21) => n_1177, data_out(20) => 
                           n_1178, data_out(19) => n_1179, data_out(18) => 
                           n_1180, data_out(17) => n_1181, data_out(16) => 
                           n_1182, data_out(15) => n_1183, data_out(14) => 
                           n_1184, data_out(13) => n_1185, data_out(12) => 
                           n_1186, data_out(11) => n_1187, data_out(10) => 
                           n_1188, data_out(9) => n_1189, data_out(8) => n_1190
                           , data_out(7) => n_1191, data_out(6) => n_1192, 
                           data_out(5) => n_1193, data_out(4) => n_1194, 
                           data_out(3) => n_1195, data_out(2) => n_1196, 
                           data_out(1) => n_1197, data_out(0) => cmp_out_0_port
                           );
   mux : mux11to1_nbit32 port map( A(31) => p4_out_31_port, A(30) => 
                           p4_out_30_port, A(29) => p4_out_29_port, A(28) => 
                           p4_out_28_port, A(27) => p4_out_27_port, A(26) => 
                           p4_out_26_port, A(25) => p4_out_25_port, A(24) => 
                           p4_out_24_port, A(23) => p4_out_23_port, A(22) => 
                           p4_out_22_port, A(21) => p4_out_21_port, A(20) => 
                           p4_out_20_port, A(19) => p4_out_19_port, A(18) => 
                           p4_out_18_port, A(17) => p4_out_17_port, A(16) => 
                           p4_out_16_port, A(15) => p4_out_15_port, A(14) => 
                           p4_out_14_port, A(13) => p4_out_13_port, A(12) => 
                           p4_out_12_port, A(11) => p4_out_11_port, A(10) => 
                           p4_out_10_port, A(9) => p4_out_9_port, A(8) => 
                           p4_out_8_port, A(7) => p4_out_7_port, A(6) => 
                           p4_out_6_port, A(5) => p4_out_5_port, A(4) => 
                           p4_out_4_port, A(3) => p4_out_3_port, A(2) => 
                           p4_out_2_port, A(1) => p4_out_1_port, A(0) => 
                           p4_out_0_port, B(31) => and_out_31_port, B(30) => 
                           and_out_30_port, B(29) => and_out_29_port, B(28) => 
                           and_out_28_port, B(27) => and_out_27_port, B(26) => 
                           and_out_26_port, B(25) => and_out_25_port, B(24) => 
                           and_out_24_port, B(23) => and_out_23_port, B(22) => 
                           and_out_22_port, B(21) => and_out_21_port, B(20) => 
                           and_out_20_port, B(19) => and_out_19_port, B(18) => 
                           and_out_18_port, B(17) => and_out_17_port, B(16) => 
                           and_out_16_port, B(15) => and_out_15_port, B(14) => 
                           and_out_14_port, B(13) => and_out_13_port, B(12) => 
                           and_out_12_port, B(11) => and_out_11_port, B(10) => 
                           and_out_10_port, B(9) => and_out_9_port, B(8) => 
                           and_out_8_port, B(7) => and_out_7_port, B(6) => 
                           and_out_6_port, B(5) => and_out_5_port, B(4) => 
                           and_out_4_port, B(3) => and_out_3_port, B(2) => 
                           and_out_2_port, B(1) => and_out_1_port, B(0) => 
                           and_out_0_port, C(31) => or_out_31_port, C(30) => 
                           or_out_30_port, C(29) => or_out_29_port, C(28) => 
                           or_out_28_port, C(27) => or_out_27_port, C(26) => 
                           or_out_26_port, C(25) => or_out_25_port, C(24) => 
                           or_out_24_port, C(23) => or_out_23_port, C(22) => 
                           or_out_22_port, C(21) => or_out_21_port, C(20) => 
                           or_out_20_port, C(19) => or_out_19_port, C(18) => 
                           or_out_18_port, C(17) => or_out_17_port, C(16) => 
                           or_out_16_port, C(15) => or_out_15_port, C(14) => 
                           or_out_14_port, C(13) => or_out_13_port, C(12) => 
                           or_out_12_port, C(11) => or_out_11_port, C(10) => 
                           or_out_10_port, C(9) => or_out_9_port, C(8) => 
                           or_out_8_port, C(7) => or_out_7_port, C(6) => 
                           or_out_6_port, C(5) => or_out_5_port, C(4) => 
                           or_out_4_port, C(3) => or_out_3_port, C(2) => 
                           or_out_2_port, C(1) => or_out_1_port, C(0) => 
                           or_out_0_port, D(31) => xor_out_31_port, D(30) => 
                           xor_out_30_port, D(29) => xor_out_29_port, D(28) => 
                           xor_out_28_port, D(27) => xor_out_27_port, D(26) => 
                           xor_out_26_port, D(25) => xor_out_25_port, D(24) => 
                           xor_out_24_port, D(23) => xor_out_23_port, D(22) => 
                           xor_out_22_port, D(21) => xor_out_21_port, D(20) => 
                           xor_out_20_port, D(19) => xor_out_19_port, D(18) => 
                           xor_out_18_port, D(17) => xor_out_17_port, D(16) => 
                           xor_out_16_port, D(15) => xor_out_15_port, D(14) => 
                           xor_out_14_port, D(13) => xor_out_13_port, D(12) => 
                           xor_out_12_port, D(11) => xor_out_11_port, D(10) => 
                           xor_out_10_port, D(9) => xor_out_9_port, D(8) => 
                           xor_out_8_port, D(7) => xor_out_7_port, D(6) => 
                           xor_out_6_port, D(5) => xor_out_5_port, D(4) => 
                           xor_out_4_port, D(3) => xor_out_3_port, D(2) => 
                           xor_out_2_port, D(1) => xor_out_1_port, D(0) => 
                           xor_out_0_port, E(31) => sl_out_31_port, E(30) => 
                           sl_out_30_port, E(29) => sl_out_29_port, E(28) => 
                           sl_out_28_port, E(27) => sl_out_27_port, E(26) => 
                           sl_out_26_port, E(25) => sl_out_25_port, E(24) => 
                           sl_out_24_port, E(23) => sl_out_23_port, E(22) => 
                           sl_out_22_port, E(21) => sl_out_21_port, E(20) => 
                           sl_out_20_port, E(19) => sl_out_19_port, E(18) => 
                           sl_out_18_port, E(17) => sl_out_17_port, E(16) => 
                           sl_out_16_port, E(15) => sl_out_15_port, E(14) => 
                           sl_out_14_port, E(13) => sl_out_13_port, E(12) => 
                           sl_out_12_port, E(11) => sl_out_11_port, E(10) => 
                           sl_out_10_port, E(9) => sl_out_9_port, E(8) => 
                           sl_out_8_port, E(7) => sl_out_7_port, E(6) => 
                           sl_out_6_port, E(5) => sl_out_5_port, E(4) => 
                           sl_out_4_port, E(3) => sl_out_3_port, E(2) => 
                           sl_out_2_port, E(1) => sl_out_1_port, E(0) => 
                           sl_out_0_port, F(31) => sr_out_31_port, F(30) => 
                           sr_out_30_port, F(29) => sr_out_29_port, F(28) => 
                           sr_out_28_port, F(27) => sr_out_27_port, F(26) => 
                           sr_out_26_port, F(25) => sr_out_25_port, F(24) => 
                           sr_out_24_port, F(23) => sr_out_23_port, F(22) => 
                           sr_out_22_port, F(21) => sr_out_21_port, F(20) => 
                           sr_out_20_port, F(19) => sr_out_19_port, F(18) => 
                           sr_out_18_port, F(17) => sr_out_17_port, F(16) => 
                           sr_out_16_port, F(15) => sr_out_15_port, F(14) => 
                           sr_out_14_port, F(13) => sr_out_13_port, F(12) => 
                           sr_out_12_port, F(11) => sr_out_11_port, F(10) => 
                           sr_out_10_port, F(9) => sr_out_9_port, F(8) => 
                           sr_out_8_port, F(7) => sr_out_7_port, F(6) => 
                           sr_out_6_port, F(5) => sr_out_5_port, F(4) => 
                           sr_out_4_port, F(3) => sr_out_3_port, F(2) => 
                           sr_out_2_port, F(1) => sr_out_1_port, F(0) => 
                           sr_out_0_port, H(31) => cmp_out_31_port, H(30) => 
                           cmp_out_30_port, H(29) => cmp_out_29_port, H(28) => 
                           cmp_out_28_port, H(27) => cmp_out_27_port, H(26) => 
                           cmp_out_26_port, H(25) => cmp_out_25_port, H(24) => 
                           cmp_out_24_port, H(23) => cmp_out_23_port, H(22) => 
                           cmp_out_22_port, H(21) => cmp_out_21_port, H(20) => 
                           cmp_out_20_port, H(19) => cmp_out_19_port, H(18) => 
                           cmp_out_18_port, H(17) => cmp_out_17_port, H(16) => 
                           cmp_out_16_port, H(15) => cmp_out_15_port, H(14) => 
                           cmp_out_14_port, H(13) => cmp_out_13_port, H(12) => 
                           cmp_out_12_port, H(11) => cmp_out_11_port, H(10) => 
                           cmp_out_10_port, H(9) => cmp_out_9_port, H(8) => 
                           cmp_out_8_port, H(7) => cmp_out_7_port, H(6) => 
                           cmp_out_6_port, H(5) => cmp_out_5_port, H(4) => 
                           cmp_out_4_port, H(3) => cmp_out_3_port, H(2) => 
                           cmp_out_2_port, H(1) => cmp_out_1_port, H(0) => 
                           cmp_out_0_port, sel(3) => mux_sel_3_port, sel(2) => 
                           mux_sel_2_port, sel(1) => mux_sel_1_port, sel(0) => 
                           mux_sel_0_port, Y(31) => data_out(31), Y(30) => 
                           data_out(30), Y(29) => data_out(29), Y(28) => 
                           data_out(28), Y(27) => data_out(27), Y(26) => 
                           data_out(26), Y(25) => data_out(25), Y(24) => 
                           data_out(24), Y(23) => data_out(23), Y(22) => 
                           data_out(22), Y(21) => data_out(21), Y(20) => 
                           data_out(20), Y(19) => data_out(19), Y(18) => 
                           data_out(18), Y(17) => data_out(17), Y(16) => 
                           data_out(16), Y(15) => data_out(15), Y(14) => 
                           data_out(14), Y(13) => data_out(13), Y(12) => 
                           data_out(12), Y(11) => data_out(11), Y(10) => 
                           data_out(10), Y(9) => data_out(9), Y(8) => 
                           data_out(8), Y(7) => data_out(7), Y(6) => 
                           data_out(6), Y(5) => data_out(5), Y(4) => 
                           data_out(4), Y(3) => data_out(3), Y(2) => 
                           data_out(2), Y(1) => data_out(1), Y(0) => 
                           data_out(0));
   add_sel_reg : DLH_X1 port map( G => N41, D => n56, Q => add_sel);
   U3 : BUF_X1 port map( A => n65, Z => n71);
   U4 : BUF_X2 port map( A => data_in2(3), Z => n63);
   U5 : BUF_X1 port map( A => data_in1(13), Z => n83);
   U6 : BUF_X1 port map( A => data_in1(14), Z => n84);
   U7 : BUF_X2 port map( A => data_in1(18), Z => n85);
   U8 : NOR4_X1 port map( A1 => n45, A2 => N49, A3 => n54, A4 => n55, ZN => n40
                           );
   U9 : BUF_X1 port map( A => data_in1(9), Z => n82);
   U10 : CLKBUF_X1 port map( A => data_in2(24), Z => n52);
   U11 : CLKBUF_X1 port map( A => data_in2(13), Z => n53);
   U12 : CLKBUF_X1 port map( A => data_in2(22), Z => n57);
   U13 : BUF_X2 port map( A => data_in2(10), Z => n58);
   U14 : CLKBUF_X1 port map( A => data_in2(7), Z => n59);
   U15 : CLKBUF_X1 port map( A => data_in2(23), Z => n60);
   U16 : BUF_X1 port map( A => data_in2(2), Z => n65);
   U17 : BUF_X2 port map( A => data_in2(30), Z => n61);
   U18 : CLKBUF_X1 port map( A => data_in2(26), Z => n62);
   U19 : CLKBUF_X1 port map( A => data_in2(28), Z => n64);
   U20 : CLKBUF_X1 port map( A => data_in1(1), Z => n66);
   U21 : CLKBUF_X1 port map( A => data_in1(0), Z => n79);
   U22 : CLKBUF_X1 port map( A => data_in2(0), Z => n72);
   U23 : INV_X1 port map( A => n69, ZN => n119);
   U24 : INV_X1 port map( A => n77, ZN => n111);
   U25 : INV_X1 port map( A => n74, ZN => n114);
   U26 : INV_X1 port map( A => n71, ZN => n118);
   U27 : INV_X1 port map( A => n73, ZN => n101);
   U28 : INV_X1 port map( A => n78, ZN => n91);
   U29 : INV_X1 port map( A => n58, ZN => n110);
   U30 : INV_X1 port map( A => n63, ZN => n117);
   U31 : INV_X1 port map( A => n62, ZN => n94);
   U32 : INV_X1 port map( A => data_in2(4), ZN => n116);
   U33 : INV_X1 port map( A => data_in2(31), ZN => n89);
   U34 : INV_X1 port map( A => data_in2(11), ZN => n109);
   U35 : INV_X1 port map( A => data_in2(12), ZN => n108);
   U36 : INV_X1 port map( A => data_in2(14), ZN => n106);
   U37 : INV_X1 port map( A => data_in2(15), ZN => n105);
   U38 : INV_X1 port map( A => n60, ZN => n97);
   U39 : INV_X1 port map( A => data_in2(17), ZN => n103);
   U40 : INV_X1 port map( A => data_in2(16), ZN => n104);
   U41 : INV_X1 port map( A => data_in2(18), ZN => n102);
   U42 : INV_X1 port map( A => data_in2(5), ZN => n115);
   U43 : INV_X1 port map( A => n61, ZN => n90);
   U44 : INV_X1 port map( A => data_in2(27), ZN => n93);
   U45 : INV_X1 port map( A => data_in2(25), ZN => n95);
   U46 : INV_X1 port map( A => data_in2(20), ZN => n100);
   U47 : INV_X1 port map( A => n59, ZN => n113);
   U48 : INV_X1 port map( A => n52, ZN => n96);
   U49 : NOR2_X1 port map( A1 => n124, A2 => n42_port, ZN => n55);
   U50 : OR3_X1 port map( A1 => n126, A2 => n127, A3 => n44_port, ZN => 
                           n43_port);
   U51 : INV_X1 port map( A => n40, ZN => n121);
   U52 : INV_X1 port map( A => n50, ZN => n122);
   U53 : NAND2_X1 port map( A1 => n41_port, A2 => n40, ZN => n50);
   U54 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => n44_port);
   U55 : INV_X1 port map( A => n41_port, ZN => n123);
   U56 : BUF_X1 port map( A => data_in1(21), Z => n86);
   U93 : BUF_X1 port map( A => data_in1(22), Z => n87);
   U94 : BUF_X1 port map( A => data_in1(30), Z => n88);
   U95 : AND2_X1 port map( A1 => n47, A2 => op_sel(1), ZN => n45);
   U96 : NOR4_X1 port map( A1 => n127, A2 => n124, A3 => n125, A4 => op_sel(1),
                           ZN => n54);
   U97 : AOI211_X1 port map( C1 => n126, C2 => n47, A => n48, B => n51, ZN => 
                           n41_port);
   U98 : NOR3_X1 port map( A1 => n125, A2 => op_sel(3), A3 => n127, ZN => n48);
   U99 : NOR3_X1 port map( A1 => op_sel(0), A2 => op_sel(2), A3 => n124, ZN => 
                           n47);
   U100 : NOR2_X1 port map( A1 => n44_port, A2 => op_sel(1), ZN => N41);
   U101 : INV_X1 port map( A => op_sel(3), ZN => n124);
   U102 : INV_X1 port map( A => op_sel(0), ZN => n127);
   U103 : INV_X1 port map( A => op_sel(2), ZN => n125);
   U104 : INV_X1 port map( A => op_sel(1), ZN => n126);
   U105 : OAI21_X1 port map( B1 => op_sel(0), B2 => N41, A => n40, ZN => N43);
   U106 : AND3_X1 port map( A1 => op_sel(3), A2 => n46, A3 => op_sel(1), ZN => 
                           N49);
   U107 : AND3_X1 port map( A1 => n49_port, A2 => n124, A3 => op_sel(2), ZN => 
                           n51);
   U108 : AND2_X1 port map( A1 => op_sel(0), A2 => N41, ZN => n56);
   U109 : CLKBUF_X1 port map( A => data_in1(2), Z => n67);
   U110 : INV_X1 port map( A => n53, ZN => n107);
   U111 : CLKBUF_X1 port map( A => data_in2(1), Z => n68);
   U112 : CLKBUF_X1 port map( A => data_in2(1), Z => n69);
   U113 : CLKBUF_X1 port map( A => n65, Z => n70);
   U114 : CLKBUF_X1 port map( A => data_in2(19), Z => n73);
   U115 : CLKBUF_X1 port map( A => data_in2(6), Z => n74);
   U116 : CLKBUF_X1 port map( A => data_in2(21), Z => n75);
   U117 : INV_X1 port map( A => n57, ZN => n98);
   U118 : CLKBUF_X1 port map( A => data_in2(8), Z => n76);
   U119 : CLKBUF_X1 port map( A => data_in2(9), Z => n77);
   U120 : CLKBUF_X1 port map( A => data_in2(29), Z => n78);
   U121 : INV_X1 port map( A => n64, ZN => n92);
   U122 : INV_X1 port map( A => n75, ZN => n99);
   U123 : INV_X1 port map( A => n72, ZN => n120);
   U124 : INV_X1 port map( A => n76, ZN => n112);
   U125 : CLKBUF_X3 port map( A => data_in1(4), Z => n80);
   U126 : CLKBUF_X3 port map( A => data_in1(8), Z => n81);

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_7 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n33, n66, n67, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n100, Z => n33);
   U2 : BUF_X1 port map( A => n100, Z => n66);
   U3 : BUF_X1 port map( A => n100, Z => n67);
   U4 : INV_X1 port map( A => n101, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n33, B1 => B(0), B2 => SEL, ZN => 
                           n101);
   U6 : INV_X1 port map( A => n112, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => n33, B1 => B(1), B2 => SEL, ZN => 
                           n112);
   U8 : INV_X1 port map( A => n119, ZN => Y(26));
   U9 : AOI22_X1 port map( A1 => A(26), A2 => n66, B1 => B(26), B2 => SEL, ZN 
                           => n119);
   U10 : INV_X1 port map( A => n120, ZN => Y(27));
   U11 : AOI22_X1 port map( A1 => A(27), A2 => n66, B1 => B(27), B2 => SEL, ZN 
                           => n120);
   U12 : INV_X1 port map( A => n121, ZN => Y(28));
   U13 : AOI22_X1 port map( A1 => A(28), A2 => n66, B1 => B(28), B2 => SEL, ZN 
                           => n121);
   U14 : INV_X1 port map( A => n122, ZN => Y(29));
   U15 : AOI22_X1 port map( A1 => A(29), A2 => n66, B1 => B(29), B2 => SEL, ZN 
                           => n122);
   U16 : INV_X1 port map( A => n124, ZN => Y(30));
   U17 : AOI22_X1 port map( A1 => A(30), A2 => n66, B1 => B(30), B2 => SEL, ZN 
                           => n124);
   U18 : INV_X1 port map( A => n125, ZN => Y(31));
   U19 : AOI22_X1 port map( A1 => A(31), A2 => n67, B1 => B(31), B2 => SEL, ZN 
                           => n125);
   U20 : INV_X1 port map( A => n104, ZN => Y(12));
   U21 : AOI22_X1 port map( A1 => A(12), A2 => n33, B1 => B(12), B2 => SEL, ZN 
                           => n104);
   U22 : INV_X1 port map( A => n105, ZN => Y(13));
   U23 : AOI22_X1 port map( A1 => A(13), A2 => n33, B1 => B(13), B2 => SEL, ZN 
                           => n105);
   U24 : INV_X1 port map( A => n106, ZN => Y(14));
   U25 : AOI22_X1 port map( A1 => A(14), A2 => n33, B1 => B(14), B2 => SEL, ZN 
                           => n106);
   U26 : INV_X1 port map( A => n107, ZN => Y(15));
   U27 : AOI22_X1 port map( A1 => A(15), A2 => n33, B1 => B(15), B2 => SEL, ZN 
                           => n107);
   U28 : INV_X1 port map( A => n108, ZN => Y(16));
   U29 : AOI22_X1 port map( A1 => A(16), A2 => n33, B1 => B(16), B2 => SEL, ZN 
                           => n108);
   U30 : INV_X1 port map( A => n109, ZN => Y(17));
   U31 : AOI22_X1 port map( A1 => A(17), A2 => n33, B1 => B(17), B2 => SEL, ZN 
                           => n109);
   U32 : INV_X1 port map( A => n110, ZN => Y(18));
   U33 : AOI22_X1 port map( A1 => A(18), A2 => n33, B1 => B(18), B2 => SEL, ZN 
                           => n110);
   U34 : INV_X1 port map( A => n111, ZN => Y(19));
   U35 : AOI22_X1 port map( A1 => A(19), A2 => n33, B1 => B(19), B2 => SEL, ZN 
                           => n111);
   U36 : INV_X1 port map( A => n113, ZN => Y(20));
   U37 : AOI22_X1 port map( A1 => A(20), A2 => n66, B1 => B(20), B2 => SEL, ZN 
                           => n113);
   U38 : INV_X1 port map( A => n114, ZN => Y(21));
   U39 : AOI22_X1 port map( A1 => A(21), A2 => n66, B1 => B(21), B2 => SEL, ZN 
                           => n114);
   U40 : INV_X1 port map( A => n115, ZN => Y(22));
   U41 : AOI22_X1 port map( A1 => A(22), A2 => n66, B1 => B(22), B2 => SEL, ZN 
                           => n115);
   U42 : INV_X1 port map( A => n116, ZN => Y(23));
   U43 : AOI22_X1 port map( A1 => A(23), A2 => n66, B1 => B(23), B2 => SEL, ZN 
                           => n116);
   U44 : INV_X1 port map( A => n117, ZN => Y(24));
   U45 : AOI22_X1 port map( A1 => A(24), A2 => n66, B1 => B(24), B2 => SEL, ZN 
                           => n117);
   U46 : INV_X1 port map( A => n118, ZN => Y(25));
   U47 : AOI22_X1 port map( A1 => A(25), A2 => n66, B1 => B(25), B2 => SEL, ZN 
                           => n118);
   U48 : INV_X1 port map( A => n123, ZN => Y(2));
   U49 : AOI22_X1 port map( A1 => A(2), A2 => n66, B1 => B(2), B2 => SEL, ZN =>
                           n123);
   U50 : INV_X1 port map( A => n126, ZN => Y(3));
   U51 : AOI22_X1 port map( A1 => A(3), A2 => n67, B1 => B(3), B2 => SEL, ZN =>
                           n126);
   U52 : INV_X1 port map( A => n127, ZN => Y(4));
   U53 : AOI22_X1 port map( A1 => A(4), A2 => n67, B1 => B(4), B2 => SEL, ZN =>
                           n127);
   U54 : INV_X1 port map( A => n128, ZN => Y(5));
   U55 : AOI22_X1 port map( A1 => A(5), A2 => n67, B1 => B(5), B2 => SEL, ZN =>
                           n128);
   U56 : INV_X1 port map( A => n129, ZN => Y(6));
   U57 : AOI22_X1 port map( A1 => A(6), A2 => n67, B1 => B(6), B2 => SEL, ZN =>
                           n129);
   U58 : INV_X1 port map( A => n130, ZN => Y(7));
   U59 : AOI22_X1 port map( A1 => A(7), A2 => n67, B1 => B(7), B2 => SEL, ZN =>
                           n130);
   U60 : INV_X1 port map( A => n131, ZN => Y(8));
   U61 : AOI22_X1 port map( A1 => A(8), A2 => n67, B1 => B(8), B2 => SEL, ZN =>
                           n131);
   U62 : INV_X1 port map( A => n132, ZN => Y(9));
   U63 : AOI22_X1 port map( A1 => A(9), A2 => n67, B1 => SEL, B2 => B(9), ZN =>
                           n132);
   U64 : INV_X1 port map( A => n102, ZN => Y(10));
   U65 : AOI22_X1 port map( A1 => A(10), A2 => n33, B1 => B(10), B2 => SEL, ZN 
                           => n102);
   U66 : INV_X1 port map( A => n103, ZN => Y(11));
   U67 : AOI22_X1 port map( A1 => A(11), A2 => n33, B1 => B(11), B2 => SEL, ZN 
                           => n103);
   U68 : INV_X1 port map( A => SEL, ZN => n100);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_8 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_8;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n33, n66, n67, n100 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n39, ZN => Y(4));
   U2 : INV_X1 port map( A => n58, ZN => Y(16));
   U3 : INV_X1 port map( A => n57, ZN => Y(17));
   U4 : INV_X1 port map( A => n56, ZN => Y(18));
   U5 : INV_X1 port map( A => n48, ZN => Y(25));
   U6 : INV_X1 port map( A => n46, ZN => Y(27));
   U7 : INV_X1 port map( A => n42, ZN => Y(30));
   U8 : INV_X1 port map( A => n64, ZN => Y(10));
   U9 : INV_X1 port map( A => n62, ZN => Y(12));
   U10 : INV_X1 port map( A => n63, ZN => Y(11));
   U11 : INV_X1 port map( A => n38, ZN => Y(5));
   U12 : INV_X1 port map( A => n40, ZN => Y(3));
   U13 : INV_X1 port map( A => n50, ZN => Y(23));
   U14 : BUF_X1 port map( A => n100, Z => n33);
   U15 : BUF_X1 port map( A => n100, Z => n66);
   U16 : BUF_X1 port map( A => n100, Z => n67);
   U17 : AOI22_X1 port map( A1 => A(3), A2 => n67, B1 => B(3), B2 => SEL, ZN =>
                           n40);
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n67, B1 => B(4), B2 => SEL, ZN =>
                           n39);
   U19 : AOI22_X1 port map( A1 => A(11), A2 => n33, B1 => B(11), B2 => SEL, ZN 
                           => n63);
   U20 : AOI22_X1 port map( A1 => A(12), A2 => n33, B1 => B(12), B2 => SEL, ZN 
                           => n62);
   U21 : AOI22_X1 port map( A1 => A(10), A2 => n33, B1 => B(10), B2 => SEL, ZN 
                           => n64);
   U22 : AOI22_X1 port map( A1 => A(17), A2 => n33, B1 => B(17), B2 => SEL, ZN 
                           => n57);
   U23 : AOI22_X1 port map( A1 => A(16), A2 => n33, B1 => B(16), B2 => SEL, ZN 
                           => n58);
   U24 : AOI22_X1 port map( A1 => A(18), A2 => n33, B1 => B(18), B2 => SEL, ZN 
                           => n56);
   U25 : AOI22_X1 port map( A1 => A(5), A2 => n67, B1 => B(5), B2 => SEL, ZN =>
                           n38);
   U26 : AOI22_X1 port map( A1 => A(30), A2 => n66, B1 => B(30), B2 => SEL, ZN 
                           => n42);
   U27 : AOI22_X1 port map( A1 => A(27), A2 => n66, B1 => B(27), B2 => SEL, ZN 
                           => n46);
   U28 : AOI22_X1 port map( A1 => A(23), A2 => n66, B1 => B(23), B2 => SEL, ZN 
                           => n50);
   U29 : AOI22_X1 port map( A1 => A(25), A2 => n66, B1 => B(25), B2 => SEL, ZN 
                           => n48);
   U30 : INV_X1 port map( A => n59, ZN => Y(15));
   U31 : AOI22_X1 port map( A1 => A(15), A2 => n33, B1 => B(15), B2 => SEL, ZN 
                           => n59);
   U32 : INV_X1 port map( A => n53, ZN => Y(20));
   U33 : AOI22_X1 port map( A1 => A(20), A2 => n66, B1 => B(20), B2 => SEL, ZN 
                           => n53);
   U34 : INV_X1 port map( A => n49, ZN => Y(24));
   U35 : AOI22_X1 port map( A1 => A(24), A2 => n66, B1 => B(24), B2 => SEL, ZN 
                           => n49);
   U36 : INV_X1 port map( A => n41, ZN => Y(31));
   U37 : AOI22_X1 port map( A1 => A(31), A2 => n67, B1 => B(31), B2 => SEL, ZN 
                           => n41);
   U38 : INV_X1 port map( A => n60, ZN => Y(14));
   U39 : AOI22_X1 port map( A1 => A(14), A2 => n33, B1 => B(14), B2 => SEL, ZN 
                           => n60);
   U40 : INV_X1 port map( A => n61, ZN => Y(13));
   U41 : AOI22_X1 port map( A1 => A(13), A2 => n33, B1 => B(13), B2 => SEL, ZN 
                           => n61);
   U42 : INV_X1 port map( A => n36, ZN => Y(7));
   U43 : AOI22_X1 port map( A1 => A(7), A2 => n67, B1 => B(7), B2 => SEL, ZN =>
                           n36);
   U44 : AOI22_X1 port map( A1 => A(9), A2 => n67, B1 => SEL, B2 => B(9), ZN =>
                           n34);
   U45 : AOI22_X1 port map( A1 => A(2), A2 => n66, B1 => B(2), B2 => SEL, ZN =>
                           n43);
   U46 : AOI22_X1 port map( A1 => A(1), A2 => n33, B1 => B(1), B2 => SEL, ZN =>
                           n54);
   U47 : AOI22_X1 port map( A1 => A(0), A2 => n33, B1 => B(0), B2 => SEL, ZN =>
                           n65);
   U48 : INV_X1 port map( A => SEL, ZN => n100);
   U49 : INV_X1 port map( A => n54, ZN => Y(1));
   U50 : INV_X1 port map( A => n43, ZN => Y(2));
   U51 : INV_X1 port map( A => n65, ZN => Y(0));
   U52 : INV_X1 port map( A => n55, ZN => Y(19));
   U53 : AOI22_X1 port map( A1 => A(26), A2 => n66, B1 => B(26), B2 => SEL, ZN 
                           => n47);
   U54 : INV_X1 port map( A => n47, ZN => Y(26));
   U55 : AOI22_X1 port map( A1 => A(19), A2 => n33, B1 => B(19), B2 => SEL, ZN 
                           => n55);
   U56 : INV_X1 port map( A => n37, ZN => Y(6));
   U57 : AOI22_X1 port map( A1 => A(6), A2 => n67, B1 => B(6), B2 => SEL, ZN =>
                           n37);
   U58 : INV_X1 port map( A => n34, ZN => Y(9));
   U59 : INV_X1 port map( A => n51, ZN => Y(22));
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n66, B1 => B(22), B2 => SEL, ZN 
                           => n51);
   U61 : INV_X1 port map( A => n44, ZN => Y(29));
   U62 : AOI22_X1 port map( A1 => A(29), A2 => n66, B1 => B(29), B2 => SEL, ZN 
                           => n44);
   U63 : AOI22_X1 port map( A1 => A(8), A2 => n67, B1 => B(8), B2 => SEL, ZN =>
                           n35);
   U64 : INV_X1 port map( A => n35, ZN => Y(8));
   U65 : INV_X1 port map( A => n45, ZN => Y(28));
   U66 : AOI22_X1 port map( A1 => A(28), A2 => n66, B1 => B(28), B2 => SEL, ZN 
                           => n45);
   U67 : AOI22_X1 port map( A1 => A(21), A2 => n66, B1 => B(21), B2 => SEL, ZN 
                           => n52);
   U68 : INV_X1 port map( A => n52, ZN => Y(21));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_10 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_10;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n50, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n50, Q => Q(30), 
                           QN => n67);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n50, Q => Q(29), 
                           QN => n68);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n50, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n50, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n50, Q => Q(26), 
                           QN => n71);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n50, Q => Q(25),
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n50, Q => Q(24),
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n50, Q => Q(23),
                           QN => n74);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n50, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n50, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n50, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n51, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n51, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n51, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n51, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n51, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n51, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n51, Q => Q(8), 
                           QN => n89);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n52, Q => Q(7), 
                           QN => n90);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n52, Q => Q(6), 
                           QN => n91);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n52, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n52, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n52, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n52, Q => Q(2), 
                           QN => n95);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n52, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n52, Q => Q(0), 
                           QN => n97);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n51);
   U5 : BUF_X1 port map( A => RESET_n, Z => n50);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n44);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n97, A2 => n40, B1 => n42, B2 => n116, ZN => 
                           n35);
   U20 : INV_X1 port map( A => D(0), ZN => n116);
   U21 : OAI22_X1 port map( A1 => n96, A2 => n39, B1 => n42, B2 => n115, ZN => 
                           n34);
   U22 : INV_X1 port map( A => D(1), ZN => n115);
   U23 : OAI22_X1 port map( A1 => n71, A2 => n40, B1 => n41, B2 => n58, ZN => 
                           n9);
   U24 : INV_X1 port map( A => D(26), ZN => n58);
   U25 : OAI22_X1 port map( A1 => n70, A2 => n39, B1 => n41, B2 => n57, ZN => 
                           n8);
   U26 : INV_X1 port map( A => D(27), ZN => n57);
   U27 : OAI22_X1 port map( A1 => n69, A2 => n40, B1 => n41, B2 => n56, ZN => 
                           n7);
   U28 : INV_X1 port map( A => D(28), ZN => n56);
   U29 : OAI22_X1 port map( A1 => n68, A2 => n39, B1 => n41, B2 => n55, ZN => 
                           n6);
   U30 : INV_X1 port map( A => D(29), ZN => n55);
   U31 : OAI22_X1 port map( A1 => n67, A2 => n40, B1 => n42, B2 => n54, ZN => 
                           n5);
   U32 : INV_X1 port map( A => D(30), ZN => n54);
   U33 : OAI22_X1 port map( A1 => n66, A2 => n39, B1 => n42, B2 => n53, ZN => 
                           n4);
   U34 : INV_X1 port map( A => D(31), ZN => n53);
   U35 : OAI22_X1 port map( A1 => n95, A2 => n40, B1 => n43, B2 => n114, ZN => 
                           n33);
   U36 : INV_X1 port map( A => D(2), ZN => n114);
   U37 : OAI22_X1 port map( A1 => n94, A2 => n40, B1 => n43, B2 => n113, ZN => 
                           n32);
   U38 : INV_X1 port map( A => D(3), ZN => n113);
   U39 : OAI22_X1 port map( A1 => n93, A2 => n40, B1 => n43, B2 => n112, ZN => 
                           n31);
   U40 : INV_X1 port map( A => D(4), ZN => n112);
   U41 : OAI22_X1 port map( A1 => n92, A2 => n40, B1 => n43, B2 => n111, ZN => 
                           n30);
   U42 : INV_X1 port map( A => D(5), ZN => n111);
   U43 : OAI22_X1 port map( A1 => n91, A2 => n40, B1 => n44, B2 => n110, ZN => 
                           n29);
   U44 : INV_X1 port map( A => D(6), ZN => n110);
   U45 : OAI22_X1 port map( A1 => n90, A2 => n40, B1 => n44, B2 => n109, ZN => 
                           n28);
   U46 : INV_X1 port map( A => D(7), ZN => n109);
   U47 : OAI22_X1 port map( A1 => n89, A2 => n40, B1 => n44, B2 => n108, ZN => 
                           n27);
   U48 : INV_X1 port map( A => D(8), ZN => n108);
   U49 : OAI22_X1 port map( A1 => n88, A2 => n40, B1 => n44, B2 => n107, ZN => 
                           n26);
   U50 : INV_X1 port map( A => D(9), ZN => n107);
   U51 : OAI22_X1 port map( A1 => n87, A2 => n40, B1 => n45, B2 => n106, ZN => 
                           n25);
   U52 : INV_X1 port map( A => D(10), ZN => n106);
   U53 : OAI22_X1 port map( A1 => n86, A2 => n40, B1 => n45, B2 => n105, ZN => 
                           n24);
   U54 : INV_X1 port map( A => D(11), ZN => n105);
   U55 : OAI22_X1 port map( A1 => n85, A2 => n40, B1 => n45, B2 => n104, ZN => 
                           n23);
   U56 : INV_X1 port map( A => D(12), ZN => n104);
   U57 : OAI22_X1 port map( A1 => n84, A2 => n40, B1 => n45, B2 => n103, ZN => 
                           n22);
   U58 : INV_X1 port map( A => D(13), ZN => n103);
   U59 : OAI22_X1 port map( A1 => n83, A2 => n39, B1 => n46, B2 => n102, ZN => 
                           n21);
   U60 : INV_X1 port map( A => D(14), ZN => n102);
   U61 : OAI22_X1 port map( A1 => n82, A2 => n39, B1 => n46, B2 => n101, ZN => 
                           n20);
   U62 : INV_X1 port map( A => D(15), ZN => n101);
   U63 : OAI22_X1 port map( A1 => n81, A2 => n39, B1 => n46, B2 => n100, ZN => 
                           n19);
   U64 : INV_X1 port map( A => D(16), ZN => n100);
   U65 : OAI22_X1 port map( A1 => n80, A2 => n39, B1 => n46, B2 => n99, ZN => 
                           n18);
   U66 : INV_X1 port map( A => D(17), ZN => n99);
   U67 : OAI22_X1 port map( A1 => n79, A2 => n39, B1 => n47, B2 => n98, ZN => 
                           n17);
   U68 : INV_X1 port map( A => D(18), ZN => n98);
   U69 : OAI22_X1 port map( A1 => n78, A2 => n39, B1 => n47, B2 => n65, ZN => 
                           n16);
   U70 : INV_X1 port map( A => D(19), ZN => n65);
   U71 : OAI22_X1 port map( A1 => n77, A2 => n39, B1 => n47, B2 => n64, ZN => 
                           n15);
   U72 : INV_X1 port map( A => D(20), ZN => n64);
   U73 : OAI22_X1 port map( A1 => n76, A2 => n39, B1 => n47, B2 => n63, ZN => 
                           n14);
   U74 : INV_X1 port map( A => D(21), ZN => n63);
   U75 : OAI22_X1 port map( A1 => n75, A2 => n39, B1 => n48, B2 => n62, ZN => 
                           n13);
   U76 : INV_X1 port map( A => D(22), ZN => n62);
   U77 : OAI22_X1 port map( A1 => n74, A2 => n39, B1 => n48, B2 => n61, ZN => 
                           n12);
   U78 : INV_X1 port map( A => D(23), ZN => n61);
   U79 : OAI22_X1 port map( A1 => n73, A2 => n39, B1 => n48, B2 => n60, ZN => 
                           n11);
   U80 : INV_X1 port map( A => D(24), ZN => n60);
   U81 : OAI22_X1 port map( A1 => n72, A2 => n39, B1 => n48, B2 => n59, ZN => 
                           n10);
   U82 : INV_X1 port map( A => D(25), ZN => n59);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_11 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_11;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_11 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n52, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n52, Q => Q(30), 
                           QN => n67);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n52, Q => Q(29), 
                           QN => n68);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n52, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n52, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n51, Q => Q(26), 
                           QN => n71);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n51, Q => Q(25),
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n51, Q => Q(24),
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n51, Q => Q(23),
                           QN => n74);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n51, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n51, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n52, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n52, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n50, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n50, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n50, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n50, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n50, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n50, Q => Q(8), 
                           QN => n89);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n50, Q => Q(7), 
                           QN => n90);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n50, Q => Q(6), 
                           QN => n91);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n50, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n50, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n50, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n50, Q => Q(2), 
                           QN => n95);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n51, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n52, Q => Q(0), 
                           QN => n97);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n50);
   U5 : BUF_X1 port map( A => RESET_n, Z => n51);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n45);
   U10 : BUF_X1 port map( A => n37, Z => n46);
   U11 : BUF_X1 port map( A => n36, Z => n42);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n37, Z => n44);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n71, A2 => n40, B1 => n41, B2 => n58, ZN => 
                           n9);
   U20 : INV_X1 port map( A => D(26), ZN => n58);
   U21 : OAI22_X1 port map( A1 => n70, A2 => n39, B1 => n41, B2 => n57, ZN => 
                           n8);
   U22 : INV_X1 port map( A => D(27), ZN => n57);
   U23 : OAI22_X1 port map( A1 => n68, A2 => n40, B1 => n41, B2 => n55, ZN => 
                           n6);
   U24 : INV_X1 port map( A => D(29), ZN => n55);
   U25 : OAI22_X1 port map( A1 => n67, A2 => n39, B1 => n42, B2 => n54, ZN => 
                           n5);
   U26 : INV_X1 port map( A => D(30), ZN => n54);
   U27 : OAI22_X1 port map( A1 => n66, A2 => n40, B1 => n42, B2 => n53, ZN => 
                           n4);
   U28 : INV_X1 port map( A => D(31), ZN => n53);
   U29 : OAI22_X1 port map( A1 => n97, A2 => n39, B1 => n42, B2 => n116, ZN => 
                           n35);
   U30 : INV_X1 port map( A => D(0), ZN => n116);
   U31 : OAI22_X1 port map( A1 => n96, A2 => n40, B1 => n42, B2 => n115, ZN => 
                           n34);
   U32 : INV_X1 port map( A => D(1), ZN => n115);
   U33 : INV_X1 port map( A => D(6), ZN => n110);
   U34 : INV_X1 port map( A => D(8), ZN => n108);
   U35 : INV_X1 port map( A => D(21), ZN => n63);
   U36 : INV_X1 port map( A => D(22), ZN => n62);
   U37 : INV_X1 port map( A => D(28), ZN => n56);
   U38 : OAI22_X1 port map( A1 => n95, A2 => n40, B1 => n43, B2 => n114, ZN => 
                           n33);
   U39 : INV_X1 port map( A => D(2), ZN => n114);
   U40 : OAI22_X1 port map( A1 => n94, A2 => n40, B1 => n43, B2 => n113, ZN => 
                           n32);
   U41 : INV_X1 port map( A => D(3), ZN => n113);
   U42 : OAI22_X1 port map( A1 => n93, A2 => n40, B1 => n43, B2 => n112, ZN => 
                           n31);
   U43 : INV_X1 port map( A => D(4), ZN => n112);
   U44 : OAI22_X1 port map( A1 => n92, A2 => n40, B1 => n43, B2 => n111, ZN => 
                           n30);
   U45 : INV_X1 port map( A => D(5), ZN => n111);
   U46 : OAI22_X1 port map( A1 => n90, A2 => n40, B1 => n44, B2 => n109, ZN => 
                           n28);
   U47 : INV_X1 port map( A => D(7), ZN => n109);
   U48 : OAI22_X1 port map( A1 => n88, A2 => n40, B1 => n44, B2 => n107, ZN => 
                           n26);
   U49 : INV_X1 port map( A => D(9), ZN => n107);
   U50 : OAI22_X1 port map( A1 => n87, A2 => n40, B1 => n45, B2 => n106, ZN => 
                           n25);
   U51 : INV_X1 port map( A => D(10), ZN => n106);
   U52 : OAI22_X1 port map( A1 => n86, A2 => n40, B1 => n45, B2 => n105, ZN => 
                           n24);
   U53 : INV_X1 port map( A => D(11), ZN => n105);
   U54 : OAI22_X1 port map( A1 => n85, A2 => n40, B1 => n45, B2 => n104, ZN => 
                           n23);
   U55 : INV_X1 port map( A => D(12), ZN => n104);
   U56 : OAI22_X1 port map( A1 => n84, A2 => n40, B1 => n45, B2 => n103, ZN => 
                           n22);
   U57 : INV_X1 port map( A => D(13), ZN => n103);
   U58 : OAI22_X1 port map( A1 => n83, A2 => n39, B1 => n46, B2 => n102, ZN => 
                           n21);
   U59 : INV_X1 port map( A => D(14), ZN => n102);
   U60 : OAI22_X1 port map( A1 => n82, A2 => n39, B1 => n46, B2 => n101, ZN => 
                           n20);
   U61 : INV_X1 port map( A => D(15), ZN => n101);
   U62 : OAI22_X1 port map( A1 => n81, A2 => n39, B1 => n46, B2 => n100, ZN => 
                           n19);
   U63 : INV_X1 port map( A => D(16), ZN => n100);
   U64 : OAI22_X1 port map( A1 => n80, A2 => n39, B1 => n46, B2 => n99, ZN => 
                           n18);
   U65 : INV_X1 port map( A => D(17), ZN => n99);
   U66 : OAI22_X1 port map( A1 => n79, A2 => n39, B1 => n47, B2 => n98, ZN => 
                           n17);
   U67 : INV_X1 port map( A => D(18), ZN => n98);
   U68 : OAI22_X1 port map( A1 => n78, A2 => n39, B1 => n47, B2 => n65, ZN => 
                           n16);
   U69 : INV_X1 port map( A => D(19), ZN => n65);
   U70 : OAI22_X1 port map( A1 => n77, A2 => n39, B1 => n47, B2 => n64, ZN => 
                           n15);
   U71 : INV_X1 port map( A => D(20), ZN => n64);
   U72 : OAI22_X1 port map( A1 => n74, A2 => n39, B1 => n48, B2 => n61, ZN => 
                           n12);
   U73 : INV_X1 port map( A => D(23), ZN => n61);
   U74 : OAI22_X1 port map( A1 => n73, A2 => n39, B1 => n48, B2 => n60, ZN => 
                           n11);
   U75 : INV_X1 port map( A => D(24), ZN => n60);
   U76 : OAI22_X1 port map( A1 => n72, A2 => n39, B1 => n48, B2 => n59, ZN => 
                           n10);
   U77 : INV_X1 port map( A => D(25), ZN => n59);
   U78 : OAI22_X1 port map( A1 => n69, A2 => n39, B1 => n41, B2 => n56, ZN => 
                           n7);
   U79 : OAI22_X1 port map( A1 => n91, A2 => n40, B1 => n44, B2 => n110, ZN => 
                           n29);
   U80 : OAI22_X1 port map( A1 => n76, A2 => n39, B1 => n47, B2 => n63, ZN => 
                           n14);
   U81 : OAI22_X1 port map( A1 => n75, A2 => n39, B1 => n48, B2 => n62, ZN => 
                           n13);
   U82 : OAI22_X1 port map( A1 => n89, A2 => n40, B1 => n44, B2 => n108, ZN => 
                           n27);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_12 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_12;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116 : 
      std_logic;

begin
   
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n52, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n52, Q => Q(18),
                           QN => n79);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n52, Q => Q(11),
                           QN => n86);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n52, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n52, Q => Q(2), 
                           QN => n95);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n51, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n51, Q => Q(21),
                           QN => n76);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n51, Q => Q(30), 
                           QN => n67);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n51, Q => Q(25),
                           QN => n72);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n50, Q => Q(13),
                           QN => n84);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n51, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n51, Q => Q(8), 
                           QN => n89);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n50, Q => Q(4), 
                           QN => n93);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n83);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n51, Q => Q(0), 
                           QN => n97);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n50, Q => Q(29), 
                           QN => n68);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n50, Q => Q(17),
                           QN => n80);
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n52, Q => Q(31), 
                           QN => n66);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n52, Q => Q(23),
                           QN => n74);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n50, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n50, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n51, Q => Q(26), 
                           QN => n71);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n52, Q => Q(24),
                           QN => n73);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n50, Q => Q(6), 
                           QN => n91);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n50, Q => Q(10),
                           QN => n87);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n50, Q => Q(7), 
                           QN => n90);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n51, Q => Q(5), 
                           QN => n92);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n82);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n50, Q => Q(1), 
                           QN => n96);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n50, Q => Q(20),
                           QN => n77);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n50, Q => Q(12),
                           QN => n85);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n50);
   U5 : BUF_X1 port map( A => RESET_n, Z => n51);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n37, Z => n44);
   U9 : BUF_X1 port map( A => n36, Z => n41);
   U10 : BUF_X1 port map( A => n37, Z => n46);
   U11 : BUF_X1 port map( A => n38, Z => n48);
   U12 : BUF_X1 port map( A => n36, Z => n42);
   U13 : BUF_X1 port map( A => n36, Z => n43);
   U14 : BUF_X1 port map( A => n37, Z => n45);
   U15 : BUF_X1 port map( A => n38, Z => n47);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n36);
   U18 : BUF_X1 port map( A => Enable_n, Z => n37);
   U19 : OAI22_X1 port map( A1 => n69, A2 => n40, B1 => n41, B2 => n56, ZN => 
                           n7);
   U20 : INV_X1 port map( A => D(28), ZN => n56);
   U21 : OAI22_X1 port map( A1 => n70, A2 => n39, B1 => n41, B2 => n57, ZN => 
                           n8);
   U22 : INV_X1 port map( A => D(27), ZN => n57);
   U23 : OAI22_X1 port map( A1 => n68, A2 => n40, B1 => n41, B2 => n55, ZN => 
                           n6);
   U24 : INV_X1 port map( A => D(29), ZN => n55);
   U25 : OAI22_X1 port map( A1 => n96, A2 => n39, B1 => n42, B2 => n115, ZN => 
                           n34);
   U26 : INV_X1 port map( A => D(1), ZN => n115);
   U27 : OAI22_X1 port map( A1 => n97, A2 => n39, B1 => n42, B2 => n116, ZN => 
                           n35);
   U28 : INV_X1 port map( A => D(0), ZN => n116);
   U29 : OAI22_X1 port map( A1 => n71, A2 => n40, B1 => n41, B2 => n58, ZN => 
                           n9);
   U30 : INV_X1 port map( A => D(26), ZN => n58);
   U31 : OAI22_X1 port map( A1 => n67, A2 => n39, B1 => n42, B2 => n54, ZN => 
                           n5);
   U32 : INV_X1 port map( A => D(30), ZN => n54);
   U33 : OAI22_X1 port map( A1 => n66, A2 => n40, B1 => n42, B2 => n53, ZN => 
                           n4);
   U34 : INV_X1 port map( A => D(31), ZN => n53);
   U35 : OAI22_X1 port map( A1 => n85, A2 => n40, B1 => n45, B2 => n104, ZN => 
                           n23);
   U36 : INV_X1 port map( A => D(12), ZN => n104);
   U37 : OAI22_X1 port map( A1 => n84, A2 => n40, B1 => n45, B2 => n103, ZN => 
                           n22);
   U38 : INV_X1 port map( A => D(13), ZN => n103);
   U39 : OAI22_X1 port map( A1 => n90, A2 => n40, B1 => n44, B2 => n109, ZN => 
                           n28);
   U40 : INV_X1 port map( A => D(7), ZN => n109);
   U41 : OAI22_X1 port map( A1 => n87, A2 => n40, B1 => n45, B2 => n106, ZN => 
                           n25);
   U42 : INV_X1 port map( A => D(10), ZN => n106);
   U43 : OAI22_X1 port map( A1 => n77, A2 => n39, B1 => n47, B2 => n64, ZN => 
                           n15);
   U44 : INV_X1 port map( A => D(20), ZN => n64);
   U45 : OAI22_X1 port map( A1 => n91, A2 => n40, B1 => n44, B2 => n110, ZN => 
                           n29);
   U46 : INV_X1 port map( A => D(6), ZN => n110);
   U47 : OAI22_X1 port map( A1 => n93, A2 => n40, B1 => n43, B2 => n112, ZN => 
                           n31);
   U48 : INV_X1 port map( A => D(4), ZN => n112);
   U49 : OAI22_X1 port map( A1 => n80, A2 => n39, B1 => n46, B2 => n99, ZN => 
                           n18);
   U50 : INV_X1 port map( A => D(17), ZN => n99);
   U51 : OAI22_X1 port map( A1 => n88, A2 => n40, B1 => n44, B2 => n107, ZN => 
                           n26);
   U52 : INV_X1 port map( A => D(9), ZN => n107);
   U53 : OAI22_X1 port map( A1 => n83, A2 => n39, B1 => n46, B2 => n102, ZN => 
                           n21);
   U54 : INV_X1 port map( A => D(14), ZN => n102);
   U55 : OAI22_X1 port map( A1 => n89, A2 => n40, B1 => n44, B2 => n108, ZN => 
                           n27);
   U56 : INV_X1 port map( A => D(8), ZN => n108);
   U57 : OAI22_X1 port map( A1 => n72, A2 => n39, B1 => n48, B2 => n59, ZN => 
                           n10);
   U58 : INV_X1 port map( A => D(25), ZN => n59);
   U59 : OAI22_X1 port map( A1 => n92, A2 => n40, B1 => n43, B2 => n111, ZN => 
                           n30);
   U60 : INV_X1 port map( A => D(5), ZN => n111);
   U61 : OAI22_X1 port map( A1 => n82, A2 => n39, B1 => n46, B2 => n101, ZN => 
                           n20);
   U62 : INV_X1 port map( A => D(15), ZN => n101);
   U63 : OAI22_X1 port map( A1 => n81, A2 => n39, B1 => n46, B2 => n100, ZN => 
                           n19);
   U64 : INV_X1 port map( A => D(16), ZN => n100);
   U65 : OAI22_X1 port map( A1 => n76, A2 => n39, B1 => n47, B2 => n63, ZN => 
                           n14);
   U66 : INV_X1 port map( A => D(21), ZN => n63);
   U67 : OAI22_X1 port map( A1 => n75, A2 => n39, B1 => n48, B2 => n62, ZN => 
                           n13);
   U68 : INV_X1 port map( A => D(22), ZN => n62);
   U69 : OAI22_X1 port map( A1 => n73, A2 => n39, B1 => n48, B2 => n60, ZN => 
                           n11);
   U70 : INV_X1 port map( A => D(24), ZN => n60);
   U71 : OAI22_X1 port map( A1 => n74, A2 => n39, B1 => n48, B2 => n61, ZN => 
                           n12);
   U72 : INV_X1 port map( A => D(23), ZN => n61);
   U73 : OAI22_X1 port map( A1 => n95, A2 => n40, B1 => n43, B2 => n114, ZN => 
                           n33);
   U74 : INV_X1 port map( A => D(2), ZN => n114);
   U75 : OAI22_X1 port map( A1 => n94, A2 => n40, B1 => n43, B2 => n113, ZN => 
                           n32);
   U76 : INV_X1 port map( A => D(3), ZN => n113);
   U77 : OAI22_X1 port map( A1 => n86, A2 => n40, B1 => n45, B2 => n105, ZN => 
                           n24);
   U78 : INV_X1 port map( A => D(11), ZN => n105);
   U79 : OAI22_X1 port map( A1 => n79, A2 => n39, B1 => n47, B2 => n98, ZN => 
                           n17);
   U80 : INV_X1 port map( A => D(18), ZN => n98);
   U81 : OAI22_X1 port map( A1 => n78, A2 => n39, B1 => n47, B2 => n65, ZN => 
                           n16);
   U82 : INV_X1 port map( A => D(19), ZN => n65);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_13 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_13;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n53, Q => Q(31), 
                           QN => n149);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n53, Q => Q(30), 
                           QN => n148);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n53, Q => Q(29), 
                           QN => n147);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n53, Q => Q(28), 
                           QN => n146);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n53, Q => Q(27), 
                           QN => n145);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n53, Q => Q(26), 
                           QN => n144);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n53, Q => Q(25),
                           QN => n143);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n53, Q => Q(24),
                           QN => n142);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n52, Q => Q(23),
                           QN => n141);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n52, Q => Q(22),
                           QN => n140);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n52, Q => Q(21),
                           QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n52, Q => Q(20),
                           QN => n138);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n52, Q => Q(19),
                           QN => n137);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n52, Q => Q(18),
                           QN => n136);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n52, Q => Q(17),
                           QN => n135);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n52, Q => Q(16),
                           QN => n134);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n52, Q => Q(15),
                           QN => n133);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n52, Q => Q(14),
                           QN => n132);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n52, Q => Q(13),
                           QN => n131);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n52, Q => Q(12),
                           QN => n130);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n51, Q => Q(11),
                           QN => n129);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n51, Q => Q(10),
                           QN => n128);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n51, Q => Q(9), 
                           QN => n127);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n51, Q => Q(8), 
                           QN => n126);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n51, Q => Q(7), 
                           QN => n125);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n51, Q => Q(6), 
                           QN => n124);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n51, Q => Q(5), 
                           QN => n123);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n51, Q => Q(4), 
                           QN => n122);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n51, Q => Q(3), 
                           QN => n121);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n51, Q => Q(2), 
                           QN => n120);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n51, Q => Q(1), 
                           QN => n119);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n51, Q => Q(0), 
                           QN => n118);
   U2 : INV_X1 port map( A => n50, ZN => n40);
   U3 : INV_X1 port map( A => n50, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n51);
   U5 : BUF_X1 port map( A => RESET_n, Z => n52);
   U6 : BUF_X1 port map( A => RESET_n, Z => n53);
   U7 : BUF_X1 port map( A => n38, Z => n50);
   U8 : BUF_X1 port map( A => n36, Z => n44);
   U9 : BUF_X1 port map( A => n37, Z => n45);
   U10 : BUF_X1 port map( A => n37, Z => n46);
   U11 : BUF_X1 port map( A => n37, Z => n47);
   U12 : BUF_X1 port map( A => n38, Z => n48);
   U13 : BUF_X1 port map( A => n38, Z => n49);
   U14 : BUF_X1 port map( A => n36, Z => n42);
   U15 : BUF_X1 port map( A => n36, Z => n43);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n144, A2 => n41, B1 => n42, B2 => n55, ZN => 
                           n9);
   U20 : INV_X1 port map( A => D(26), ZN => n55);
   U21 : OAI22_X1 port map( A1 => n145, A2 => n41, B1 => n42, B2 => n56, ZN => 
                           n8);
   U22 : INV_X1 port map( A => D(27), ZN => n56);
   U23 : OAI22_X1 port map( A1 => n146, A2 => n41, B1 => n42, B2 => n57, ZN => 
                           n7);
   U24 : INV_X1 port map( A => D(28), ZN => n57);
   U25 : OAI22_X1 port map( A1 => n147, A2 => n41, B1 => n42, B2 => n58, ZN => 
                           n6);
   U26 : INV_X1 port map( A => D(29), ZN => n58);
   U27 : OAI22_X1 port map( A1 => n148, A2 => n41, B1 => n43, B2 => n59, ZN => 
                           n5);
   U28 : INV_X1 port map( A => D(30), ZN => n59);
   U29 : OAI22_X1 port map( A1 => n149, A2 => n41, B1 => n43, B2 => n60, ZN => 
                           n4);
   U30 : INV_X1 port map( A => D(31), ZN => n60);
   U31 : OAI22_X1 port map( A1 => n119, A2 => n41, B1 => n43, B2 => n116, ZN =>
                           n34);
   U32 : INV_X1 port map( A => D(1), ZN => n116);
   U33 : OAI22_X1 port map( A1 => n118, A2 => n41, B1 => n43, B2 => n117, ZN =>
                           n35);
   U34 : INV_X1 port map( A => D(0), ZN => n117);
   U35 : OAI22_X1 port map( A1 => n133, A2 => n39, B1 => n47, B2 => n102, ZN =>
                           n20);
   U36 : INV_X1 port map( A => D(15), ZN => n102);
   U37 : OAI22_X1 port map( A1 => n143, A2 => n39, B1 => n49, B2 => n54, ZN => 
                           n10);
   U38 : INV_X1 port map( A => D(25), ZN => n54);
   U39 : OAI22_X1 port map( A1 => n122, A2 => n40, B1 => n44, B2 => n113, ZN =>
                           n31);
   U40 : INV_X1 port map( A => D(4), ZN => n113);
   U41 : OAI22_X1 port map( A1 => n126, A2 => n40, B1 => n45, B2 => n109, ZN =>
                           n27);
   U42 : INV_X1 port map( A => D(8), ZN => n109);
   U43 : OAI22_X1 port map( A1 => n127, A2 => n40, B1 => n45, B2 => n108, ZN =>
                           n26);
   U44 : INV_X1 port map( A => D(9), ZN => n108);
   U45 : OAI22_X1 port map( A1 => n128, A2 => n40, B1 => n46, B2 => n107, ZN =>
                           n25);
   U46 : INV_X1 port map( A => D(10), ZN => n107);
   U47 : OAI22_X1 port map( A1 => n129, A2 => n40, B1 => n46, B2 => n106, ZN =>
                           n24);
   U48 : INV_X1 port map( A => D(11), ZN => n106);
   U49 : OAI22_X1 port map( A1 => n130, A2 => n40, B1 => n46, B2 => n105, ZN =>
                           n23);
   U50 : INV_X1 port map( A => D(12), ZN => n105);
   U51 : OAI22_X1 port map( A1 => n131, A2 => n40, B1 => n46, B2 => n104, ZN =>
                           n22);
   U52 : INV_X1 port map( A => D(13), ZN => n104);
   U53 : OAI22_X1 port map( A1 => n132, A2 => n39, B1 => n47, B2 => n103, ZN =>
                           n21);
   U54 : INV_X1 port map( A => D(14), ZN => n103);
   U55 : OAI22_X1 port map( A1 => n120, A2 => n40, B1 => n44, B2 => n115, ZN =>
                           n33);
   U56 : INV_X1 port map( A => D(2), ZN => n115);
   U57 : OAI22_X1 port map( A1 => n121, A2 => n40, B1 => n44, B2 => n114, ZN =>
                           n32);
   U58 : INV_X1 port map( A => D(3), ZN => n114);
   U59 : OAI22_X1 port map( A1 => n123, A2 => n40, B1 => n44, B2 => n112, ZN =>
                           n30);
   U60 : INV_X1 port map( A => D(5), ZN => n112);
   U61 : OAI22_X1 port map( A1 => n124, A2 => n40, B1 => n45, B2 => n111, ZN =>
                           n29);
   U62 : INV_X1 port map( A => D(6), ZN => n111);
   U63 : OAI22_X1 port map( A1 => n125, A2 => n40, B1 => n45, B2 => n110, ZN =>
                           n28);
   U64 : INV_X1 port map( A => D(7), ZN => n110);
   U65 : OAI22_X1 port map( A1 => n134, A2 => n39, B1 => n47, B2 => n101, ZN =>
                           n19);
   U66 : INV_X1 port map( A => D(16), ZN => n101);
   U67 : OAI22_X1 port map( A1 => n135, A2 => n39, B1 => n47, B2 => n100, ZN =>
                           n18);
   U68 : INV_X1 port map( A => D(17), ZN => n100);
   U69 : OAI22_X1 port map( A1 => n136, A2 => n39, B1 => n48, B2 => n99, ZN => 
                           n17);
   U70 : INV_X1 port map( A => D(18), ZN => n99);
   U71 : OAI22_X1 port map( A1 => n137, A2 => n39, B1 => n48, B2 => n98, ZN => 
                           n16);
   U72 : INV_X1 port map( A => D(19), ZN => n98);
   U73 : OAI22_X1 port map( A1 => n139, A2 => n39, B1 => n48, B2 => n64, ZN => 
                           n14);
   U74 : INV_X1 port map( A => D(21), ZN => n64);
   U75 : OAI22_X1 port map( A1 => n140, A2 => n39, B1 => n49, B2 => n63, ZN => 
                           n13);
   U76 : INV_X1 port map( A => D(22), ZN => n63);
   U77 : OAI22_X1 port map( A1 => n141, A2 => n39, B1 => n49, B2 => n62, ZN => 
                           n12);
   U78 : INV_X1 port map( A => D(23), ZN => n62);
   U79 : OAI22_X1 port map( A1 => n142, A2 => n39, B1 => n49, B2 => n61, ZN => 
                           n11);
   U80 : INV_X1 port map( A => D(24), ZN => n61);
   U81 : OAI22_X1 port map( A1 => n138, A2 => n39, B1 => n48, B2 => n65, ZN => 
                           n15);
   U82 : INV_X1 port map( A => D(20), ZN => n65);
   U83 : INV_X1 port map( A => n50, ZN => n41);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_14 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_14;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n51, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n51, Q => Q(30), 
                           QN => n67);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n51, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n51, Q => Q(27), 
                           QN => n70);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n51, Q => Q(25),
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n51, Q => Q(24),
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n51, Q => Q(23),
                           QN => n74);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n52, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n52, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n52, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n52, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n52, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n52, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n52, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n51, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n51, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n50, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n50, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n50, Q => Q(9), 
                           QN => n88);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n50, Q => Q(7), 
                           QN => n90);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n50, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n50, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n50, Q => Q(3), 
                           QN => n94);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n50, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n50, Q => Q(0), 
                           QN => n97);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n51, Q => Q(29), 
                           QN => n68);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n50, Q => Q(6), 
                           QN => n91);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n51, Q => Q(26), 
                           QN => n71);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n52, Q => Q(22),
                           QN => n75);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n50, Q => Q(8), 
                           QN => n89);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n50, Q => Q(2), 
                           QN => n95);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n51);
   U5 : BUF_X1 port map( A => RESET_n, Z => n50);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n37, Z => n44);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n38, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n36, Z => n41);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n37);
   U18 : BUF_X1 port map( A => Enable_n, Z => n36);
   U19 : OAI22_X1 port map( A1 => n71, A2 => n40, B1 => n41, B2 => n64, ZN => 
                           n9);
   U20 : INV_X1 port map( A => D(26), ZN => n64);
   U21 : OAI22_X1 port map( A1 => n68, A2 => n39, B1 => n41, B2 => n99, ZN => 
                           n6);
   U22 : INV_X1 port map( A => D(29), ZN => n99);
   U23 : OAI22_X1 port map( A1 => n70, A2 => n40, B1 => n41, B2 => n65, ZN => 
                           n8);
   U24 : INV_X1 port map( A => D(27), ZN => n65);
   U25 : OAI22_X1 port map( A1 => n69, A2 => n39, B1 => n41, B2 => n98, ZN => 
                           n7);
   U26 : INV_X1 port map( A => D(28), ZN => n98);
   U27 : OAI22_X1 port map( A1 => n67, A2 => n40, B1 => n42, B2 => n100, ZN => 
                           n5);
   U28 : INV_X1 port map( A => D(30), ZN => n100);
   U29 : OAI22_X1 port map( A1 => n66, A2 => n39, B1 => n42, B2 => n101, ZN => 
                           n4);
   U30 : INV_X1 port map( A => D(31), ZN => n101);
   U31 : OAI22_X1 port map( A1 => n96, A2 => n40, B1 => n42, B2 => n115, ZN => 
                           n34);
   U32 : INV_X1 port map( A => D(1), ZN => n115);
   U33 : OAI22_X1 port map( A1 => n97, A2 => n39, B1 => n42, B2 => n116, ZN => 
                           n35);
   U34 : INV_X1 port map( A => D(0), ZN => n116);
   U35 : OAI22_X1 port map( A1 => n82, A2 => n39, B1 => n46, B2 => n53, ZN => 
                           n20);
   U36 : INV_X1 port map( A => D(15), ZN => n53);
   U37 : OAI22_X1 port map( A1 => n81, A2 => n39, B1 => n46, B2 => n54, ZN => 
                           n19);
   U38 : INV_X1 port map( A => D(16), ZN => n54);
   U39 : OAI22_X1 port map( A1 => n80, A2 => n39, B1 => n46, B2 => n55, ZN => 
                           n18);
   U40 : INV_X1 port map( A => D(17), ZN => n55);
   U41 : OAI22_X1 port map( A1 => n79, A2 => n39, B1 => n47, B2 => n56, ZN => 
                           n17);
   U42 : INV_X1 port map( A => D(18), ZN => n56);
   U43 : OAI22_X1 port map( A1 => n78, A2 => n39, B1 => n47, B2 => n57, ZN => 
                           n16);
   U44 : INV_X1 port map( A => D(19), ZN => n57);
   U45 : OAI22_X1 port map( A1 => n77, A2 => n39, B1 => n47, B2 => n58, ZN => 
                           n15);
   U46 : INV_X1 port map( A => D(20), ZN => n58);
   U47 : OAI22_X1 port map( A1 => n76, A2 => n39, B1 => n47, B2 => n59, ZN => 
                           n14);
   U48 : INV_X1 port map( A => D(21), ZN => n59);
   U49 : OAI22_X1 port map( A1 => n75, A2 => n39, B1 => n48, B2 => n60, ZN => 
                           n13);
   U50 : INV_X1 port map( A => D(22), ZN => n60);
   U51 : OAI22_X1 port map( A1 => n74, A2 => n39, B1 => n48, B2 => n61, ZN => 
                           n12);
   U52 : INV_X1 port map( A => D(23), ZN => n61);
   U53 : OAI22_X1 port map( A1 => n73, A2 => n39, B1 => n48, B2 => n62, ZN => 
                           n11);
   U54 : INV_X1 port map( A => D(24), ZN => n62);
   U55 : OAI22_X1 port map( A1 => n72, A2 => n39, B1 => n48, B2 => n63, ZN => 
                           n10);
   U56 : INV_X1 port map( A => D(25), ZN => n63);
   U57 : OAI22_X1 port map( A1 => n91, A2 => n40, B1 => n44, B2 => n110, ZN => 
                           n29);
   U58 : INV_X1 port map( A => D(6), ZN => n110);
   U59 : OAI22_X1 port map( A1 => n90, A2 => n40, B1 => n44, B2 => n109, ZN => 
                           n28);
   U60 : INV_X1 port map( A => D(7), ZN => n109);
   U61 : OAI22_X1 port map( A1 => n89, A2 => n40, B1 => n44, B2 => n108, ZN => 
                           n27);
   U62 : INV_X1 port map( A => D(8), ZN => n108);
   U63 : OAI22_X1 port map( A1 => n88, A2 => n40, B1 => n44, B2 => n107, ZN => 
                           n26);
   U64 : INV_X1 port map( A => D(9), ZN => n107);
   U65 : OAI22_X1 port map( A1 => n87, A2 => n40, B1 => n45, B2 => n106, ZN => 
                           n25);
   U66 : INV_X1 port map( A => D(10), ZN => n106);
   U67 : OAI22_X1 port map( A1 => n86, A2 => n40, B1 => n45, B2 => n105, ZN => 
                           n24);
   U68 : INV_X1 port map( A => D(11), ZN => n105);
   U69 : OAI22_X1 port map( A1 => n85, A2 => n40, B1 => n45, B2 => n104, ZN => 
                           n23);
   U70 : INV_X1 port map( A => D(12), ZN => n104);
   U71 : OAI22_X1 port map( A1 => n84, A2 => n40, B1 => n45, B2 => n103, ZN => 
                           n22);
   U72 : INV_X1 port map( A => D(13), ZN => n103);
   U73 : OAI22_X1 port map( A1 => n83, A2 => n39, B1 => n46, B2 => n102, ZN => 
                           n21);
   U74 : INV_X1 port map( A => D(14), ZN => n102);
   U75 : OAI22_X1 port map( A1 => n94, A2 => n40, B1 => n43, B2 => n113, ZN => 
                           n32);
   U76 : INV_X1 port map( A => D(3), ZN => n113);
   U77 : OAI22_X1 port map( A1 => n93, A2 => n40, B1 => n43, B2 => n112, ZN => 
                           n31);
   U78 : INV_X1 port map( A => D(4), ZN => n112);
   U79 : OAI22_X1 port map( A1 => n95, A2 => n40, B1 => n43, B2 => n114, ZN => 
                           n33);
   U80 : INV_X1 port map( A => D(2), ZN => n114);
   U81 : OAI22_X1 port map( A1 => n92, A2 => n40, B1 => n43, B2 => n111, ZN => 
                           n30);
   U82 : INV_X1 port map( A => D(5), ZN => n111);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_15 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_15;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n53, Q => Q(31), 
                           QN => n149);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n53, Q => Q(30), 
                           QN => n148);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n53, Q => Q(29), 
                           QN => n147);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n53, Q => Q(28), 
                           QN => n146);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n53, Q => Q(27), 
                           QN => n145);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n53, Q => Q(26), 
                           QN => n144);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n53, Q => Q(25),
                           QN => n143);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n53, Q => Q(24),
                           QN => n142);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n52, Q => Q(23),
                           QN => n141);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n52, Q => Q(22),
                           QN => n140);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n52, Q => Q(21),
                           QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n52, Q => Q(20),
                           QN => n138);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n52, Q => Q(19),
                           QN => n137);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n52, Q => Q(18),
                           QN => n136);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n52, Q => Q(17),
                           QN => n135);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n52, Q => Q(16),
                           QN => n134);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n52, Q => Q(15),
                           QN => n133);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n52, Q => Q(14),
                           QN => n132);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n52, Q => Q(13),
                           QN => n131);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n52, Q => Q(12),
                           QN => n130);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n51, Q => Q(11),
                           QN => n129);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n51, Q => Q(10),
                           QN => n128);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n51, Q => Q(9), 
                           QN => n127);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n51, Q => Q(8), 
                           QN => n126);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n51, Q => Q(7), 
                           QN => n125);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n51, Q => Q(6), 
                           QN => n124);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n51, Q => Q(5), 
                           QN => n123);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n51, Q => Q(4), 
                           QN => n122);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n51, Q => Q(3), 
                           QN => n121);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n51, Q => Q(2), 
                           QN => n120);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n51, Q => Q(1), 
                           QN => n119);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n51, Q => Q(0), 
                           QN => n118);
   U2 : INV_X1 port map( A => n50, ZN => n40);
   U3 : INV_X1 port map( A => n50, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n51);
   U5 : BUF_X1 port map( A => RESET_n, Z => n52);
   U6 : BUF_X1 port map( A => RESET_n, Z => n53);
   U7 : BUF_X1 port map( A => n38, Z => n50);
   U8 : BUF_X1 port map( A => n36, Z => n44);
   U9 : BUF_X1 port map( A => n36, Z => n43);
   U10 : BUF_X1 port map( A => n37, Z => n45);
   U11 : BUF_X1 port map( A => n37, Z => n46);
   U12 : BUF_X1 port map( A => n37, Z => n47);
   U13 : BUF_X1 port map( A => n38, Z => n48);
   U14 : BUF_X1 port map( A => n38, Z => n49);
   U15 : BUF_X1 port map( A => n36, Z => n42);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n36);
   U18 : BUF_X1 port map( A => Enable_n, Z => n37);
   U19 : OAI22_X1 port map( A1 => n118, A2 => n41, B1 => n43, B2 => n58, ZN => 
                           n35);
   U20 : INV_X1 port map( A => D(0), ZN => n58);
   U21 : OAI22_X1 port map( A1 => n119, A2 => n41, B1 => n43, B2 => n57, ZN => 
                           n34);
   U22 : INV_X1 port map( A => D(1), ZN => n57);
   U23 : OAI22_X1 port map( A1 => n144, A2 => n41, B1 => n42, B2 => n112, ZN =>
                           n9);
   U24 : INV_X1 port map( A => D(26), ZN => n112);
   U25 : OAI22_X1 port map( A1 => n145, A2 => n41, B1 => n42, B2 => n113, ZN =>
                           n8);
   U26 : INV_X1 port map( A => D(27), ZN => n113);
   U27 : OAI22_X1 port map( A1 => n146, A2 => n41, B1 => n42, B2 => n114, ZN =>
                           n7);
   U28 : INV_X1 port map( A => D(28), ZN => n114);
   U29 : OAI22_X1 port map( A1 => n147, A2 => n41, B1 => n42, B2 => n115, ZN =>
                           n6);
   U30 : INV_X1 port map( A => D(29), ZN => n115);
   U31 : OAI22_X1 port map( A1 => n148, A2 => n41, B1 => n43, B2 => n116, ZN =>
                           n5);
   U32 : INV_X1 port map( A => D(30), ZN => n116);
   U33 : OAI22_X1 port map( A1 => n149, A2 => n41, B1 => n43, B2 => n117, ZN =>
                           n4);
   U34 : INV_X1 port map( A => D(31), ZN => n117);
   U35 : OAI22_X1 port map( A1 => n120, A2 => n40, B1 => n44, B2 => n56, ZN => 
                           n33);
   U36 : INV_X1 port map( A => D(2), ZN => n56);
   U37 : OAI22_X1 port map( A1 => n121, A2 => n40, B1 => n44, B2 => n55, ZN => 
                           n32);
   U38 : INV_X1 port map( A => D(3), ZN => n55);
   U39 : OAI22_X1 port map( A1 => n122, A2 => n40, B1 => n44, B2 => n54, ZN => 
                           n31);
   U40 : INV_X1 port map( A => D(4), ZN => n54);
   U41 : OAI22_X1 port map( A1 => n123, A2 => n40, B1 => n44, B2 => n59, ZN => 
                           n30);
   U42 : INV_X1 port map( A => D(5), ZN => n59);
   U43 : OAI22_X1 port map( A1 => n124, A2 => n40, B1 => n45, B2 => n60, ZN => 
                           n29);
   U44 : INV_X1 port map( A => D(6), ZN => n60);
   U45 : OAI22_X1 port map( A1 => n125, A2 => n40, B1 => n45, B2 => n61, ZN => 
                           n28);
   U46 : INV_X1 port map( A => D(7), ZN => n61);
   U47 : OAI22_X1 port map( A1 => n126, A2 => n40, B1 => n45, B2 => n62, ZN => 
                           n27);
   U48 : INV_X1 port map( A => D(8), ZN => n62);
   U49 : OAI22_X1 port map( A1 => n127, A2 => n40, B1 => n45, B2 => n63, ZN => 
                           n26);
   U50 : INV_X1 port map( A => D(9), ZN => n63);
   U51 : OAI22_X1 port map( A1 => n128, A2 => n40, B1 => n46, B2 => n64, ZN => 
                           n25);
   U52 : INV_X1 port map( A => D(10), ZN => n64);
   U53 : OAI22_X1 port map( A1 => n129, A2 => n40, B1 => n46, B2 => n65, ZN => 
                           n24);
   U54 : INV_X1 port map( A => D(11), ZN => n65);
   U55 : OAI22_X1 port map( A1 => n130, A2 => n40, B1 => n46, B2 => n98, ZN => 
                           n23);
   U56 : INV_X1 port map( A => D(12), ZN => n98);
   U57 : OAI22_X1 port map( A1 => n131, A2 => n40, B1 => n46, B2 => n99, ZN => 
                           n22);
   U58 : INV_X1 port map( A => D(13), ZN => n99);
   U59 : OAI22_X1 port map( A1 => n132, A2 => n39, B1 => n47, B2 => n100, ZN =>
                           n21);
   U60 : INV_X1 port map( A => D(14), ZN => n100);
   U61 : OAI22_X1 port map( A1 => n133, A2 => n39, B1 => n47, B2 => n101, ZN =>
                           n20);
   U62 : INV_X1 port map( A => D(15), ZN => n101);
   U63 : OAI22_X1 port map( A1 => n134, A2 => n39, B1 => n47, B2 => n102, ZN =>
                           n19);
   U64 : INV_X1 port map( A => D(16), ZN => n102);
   U65 : OAI22_X1 port map( A1 => n135, A2 => n39, B1 => n47, B2 => n103, ZN =>
                           n18);
   U66 : INV_X1 port map( A => D(17), ZN => n103);
   U67 : OAI22_X1 port map( A1 => n136, A2 => n39, B1 => n48, B2 => n104, ZN =>
                           n17);
   U68 : INV_X1 port map( A => D(18), ZN => n104);
   U69 : OAI22_X1 port map( A1 => n137, A2 => n39, B1 => n48, B2 => n105, ZN =>
                           n16);
   U70 : INV_X1 port map( A => D(19), ZN => n105);
   U71 : OAI22_X1 port map( A1 => n138, A2 => n39, B1 => n48, B2 => n106, ZN =>
                           n15);
   U72 : INV_X1 port map( A => D(20), ZN => n106);
   U73 : OAI22_X1 port map( A1 => n139, A2 => n39, B1 => n48, B2 => n107, ZN =>
                           n14);
   U74 : INV_X1 port map( A => D(21), ZN => n107);
   U75 : OAI22_X1 port map( A1 => n140, A2 => n39, B1 => n49, B2 => n108, ZN =>
                           n13);
   U76 : INV_X1 port map( A => D(22), ZN => n108);
   U77 : OAI22_X1 port map( A1 => n141, A2 => n39, B1 => n49, B2 => n109, ZN =>
                           n12);
   U78 : INV_X1 port map( A => D(23), ZN => n109);
   U79 : OAI22_X1 port map( A1 => n142, A2 => n39, B1 => n49, B2 => n110, ZN =>
                           n11);
   U80 : INV_X1 port map( A => D(24), ZN => n110);
   U81 : OAI22_X1 port map( A1 => n143, A2 => n39, B1 => n49, B2 => n111, ZN =>
                           n10);
   U82 : INV_X1 port map( A => D(25), ZN => n111);
   U83 : INV_X1 port map( A => n50, ZN => n41);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_16 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_16;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n52, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n52, Q => Q(30), 
                           QN => n67);
   Q_reg_29_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n52, Q => Q(29), 
                           QN => n68);
   Q_reg_28_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n52, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n52, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n52, Q => Q(26), 
                           QN => n71);
   Q_reg_25_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n52, Q => Q(25),
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n52, Q => Q(24),
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n51, Q => Q(23),
                           QN => n74);
   Q_reg_22_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n51, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n51, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n51, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n51, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n51, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n51, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n51, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n51, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n51, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n51, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n51, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n50, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n50, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n50, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n50, Q => Q(8), 
                           QN => n89);
   Q_reg_7_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n50, Q => Q(7), 
                           QN => n90);
   Q_reg_6_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n50, Q => Q(6), 
                           QN => n91);
   Q_reg_5_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n50, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n50, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n50, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n33, CK => CK, RN => n50, Q => Q(2), 
                           QN => n95);
   Q_reg_1_inst : DFFR_X1 port map( D => n34, CK => CK, RN => n50, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => CK, RN => n50, Q => Q(0), 
                           QN => n97);
   U2 : INV_X1 port map( A => n49, ZN => n40);
   U3 : INV_X1 port map( A => n49, ZN => n39);
   U4 : BUF_X1 port map( A => RESET_n, Z => n50);
   U5 : BUF_X1 port map( A => RESET_n, Z => n51);
   U6 : BUF_X1 port map( A => RESET_n, Z => n52);
   U7 : BUF_X1 port map( A => n38, Z => n49);
   U8 : BUF_X1 port map( A => n36, Z => n43);
   U9 : BUF_X1 port map( A => n36, Z => n42);
   U10 : BUF_X1 port map( A => n37, Z => n44);
   U11 : BUF_X1 port map( A => n37, Z => n45);
   U12 : BUF_X1 port map( A => n37, Z => n46);
   U13 : BUF_X1 port map( A => n38, Z => n47);
   U14 : BUF_X1 port map( A => n38, Z => n48);
   U15 : BUF_X1 port map( A => n36, Z => n41);
   U16 : BUF_X1 port map( A => Enable_n, Z => n38);
   U17 : BUF_X1 port map( A => Enable_n, Z => n36);
   U18 : BUF_X1 port map( A => Enable_n, Z => n37);
   U19 : OAI22_X1 port map( A1 => n97, A2 => n39, B1 => n42, B2 => n57, ZN => 
                           n35);
   U20 : INV_X1 port map( A => D(0), ZN => n57);
   U21 : OAI22_X1 port map( A1 => n96, A2 => n40, B1 => n42, B2 => n56, ZN => 
                           n34);
   U22 : INV_X1 port map( A => D(1), ZN => n56);
   U23 : OAI22_X1 port map( A1 => n71, A2 => n40, B1 => n41, B2 => n111, ZN => 
                           n9);
   U24 : INV_X1 port map( A => D(26), ZN => n111);
   U25 : OAI22_X1 port map( A1 => n70, A2 => n39, B1 => n41, B2 => n112, ZN => 
                           n8);
   U26 : INV_X1 port map( A => D(27), ZN => n112);
   U27 : OAI22_X1 port map( A1 => n69, A2 => n40, B1 => n41, B2 => n113, ZN => 
                           n7);
   U28 : INV_X1 port map( A => D(28), ZN => n113);
   U29 : OAI22_X1 port map( A1 => n68, A2 => n39, B1 => n41, B2 => n114, ZN => 
                           n6);
   U30 : INV_X1 port map( A => D(29), ZN => n114);
   U31 : OAI22_X1 port map( A1 => n67, A2 => n40, B1 => n42, B2 => n115, ZN => 
                           n5);
   U32 : INV_X1 port map( A => D(30), ZN => n115);
   U33 : OAI22_X1 port map( A1 => n66, A2 => n39, B1 => n42, B2 => n116, ZN => 
                           n4);
   U34 : INV_X1 port map( A => D(31), ZN => n116);
   U35 : OAI22_X1 port map( A1 => n93, A2 => n40, B1 => n43, B2 => n53, ZN => 
                           n31);
   U36 : INV_X1 port map( A => D(4), ZN => n53);
   U37 : OAI22_X1 port map( A1 => n95, A2 => n40, B1 => n43, B2 => n55, ZN => 
                           n33);
   U38 : INV_X1 port map( A => D(2), ZN => n55);
   U39 : OAI22_X1 port map( A1 => n94, A2 => n40, B1 => n43, B2 => n54, ZN => 
                           n32);
   U40 : INV_X1 port map( A => D(3), ZN => n54);
   U41 : OAI22_X1 port map( A1 => n92, A2 => n40, B1 => n43, B2 => n58, ZN => 
                           n30);
   U42 : INV_X1 port map( A => D(5), ZN => n58);
   U43 : OAI22_X1 port map( A1 => n91, A2 => n40, B1 => n44, B2 => n59, ZN => 
                           n29);
   U44 : INV_X1 port map( A => D(6), ZN => n59);
   U45 : OAI22_X1 port map( A1 => n90, A2 => n40, B1 => n44, B2 => n60, ZN => 
                           n28);
   U46 : INV_X1 port map( A => D(7), ZN => n60);
   U47 : OAI22_X1 port map( A1 => n89, A2 => n40, B1 => n44, B2 => n61, ZN => 
                           n27);
   U48 : INV_X1 port map( A => D(8), ZN => n61);
   U49 : OAI22_X1 port map( A1 => n88, A2 => n40, B1 => n44, B2 => n62, ZN => 
                           n26);
   U50 : INV_X1 port map( A => D(9), ZN => n62);
   U51 : OAI22_X1 port map( A1 => n87, A2 => n40, B1 => n45, B2 => n63, ZN => 
                           n25);
   U52 : INV_X1 port map( A => D(10), ZN => n63);
   U53 : OAI22_X1 port map( A1 => n86, A2 => n40, B1 => n45, B2 => n64, ZN => 
                           n24);
   U54 : INV_X1 port map( A => D(11), ZN => n64);
   U55 : OAI22_X1 port map( A1 => n85, A2 => n40, B1 => n45, B2 => n65, ZN => 
                           n23);
   U56 : INV_X1 port map( A => D(12), ZN => n65);
   U57 : OAI22_X1 port map( A1 => n84, A2 => n40, B1 => n45, B2 => n98, ZN => 
                           n22);
   U58 : INV_X1 port map( A => D(13), ZN => n98);
   U59 : OAI22_X1 port map( A1 => n83, A2 => n39, B1 => n46, B2 => n99, ZN => 
                           n21);
   U60 : INV_X1 port map( A => D(14), ZN => n99);
   U61 : OAI22_X1 port map( A1 => n82, A2 => n39, B1 => n46, B2 => n100, ZN => 
                           n20);
   U62 : INV_X1 port map( A => D(15), ZN => n100);
   U63 : OAI22_X1 port map( A1 => n81, A2 => n39, B1 => n46, B2 => n101, ZN => 
                           n19);
   U64 : INV_X1 port map( A => D(16), ZN => n101);
   U65 : OAI22_X1 port map( A1 => n80, A2 => n39, B1 => n46, B2 => n102, ZN => 
                           n18);
   U66 : INV_X1 port map( A => D(17), ZN => n102);
   U67 : OAI22_X1 port map( A1 => n79, A2 => n39, B1 => n47, B2 => n103, ZN => 
                           n17);
   U68 : INV_X1 port map( A => D(18), ZN => n103);
   U69 : OAI22_X1 port map( A1 => n78, A2 => n39, B1 => n47, B2 => n104, ZN => 
                           n16);
   U70 : INV_X1 port map( A => D(19), ZN => n104);
   U71 : OAI22_X1 port map( A1 => n77, A2 => n39, B1 => n47, B2 => n105, ZN => 
                           n15);
   U72 : INV_X1 port map( A => D(20), ZN => n105);
   U73 : OAI22_X1 port map( A1 => n76, A2 => n39, B1 => n47, B2 => n106, ZN => 
                           n14);
   U74 : INV_X1 port map( A => D(21), ZN => n106);
   U75 : OAI22_X1 port map( A1 => n75, A2 => n39, B1 => n48, B2 => n107, ZN => 
                           n13);
   U76 : INV_X1 port map( A => D(22), ZN => n107);
   U77 : OAI22_X1 port map( A1 => n74, A2 => n39, B1 => n48, B2 => n108, ZN => 
                           n12);
   U78 : INV_X1 port map( A => D(23), ZN => n108);
   U79 : OAI22_X1 port map( A1 => n73, A2 => n39, B1 => n48, B2 => n109, ZN => 
                           n11);
   U80 : INV_X1 port map( A => D(24), ZN => n109);
   U81 : OAI22_X1 port map( A1 => n72, A2 => n39, B1 => n48, B2 => n110, ZN => 
                           n10);
   U82 : INV_X1 port map( A => D(25), ZN => n110);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity sign_extension_sign_init16_sign_ext32 is

   port( data_in : in std_logic_vector (15 downto 0);  data_out : out 
         std_logic_vector (31 downto 0));

end sign_extension_sign_init16_sign_ext32;

architecture SYN_BEH of sign_extension_sign_init16_sign_ext32 is

begin
   data_out <= ( data_in(15), data_in(15), data_in(15), data_in(15), 
      data_in(15), data_in(15), data_in(15), data_in(15), data_in(15), 
      data_in(15), data_in(15), data_in(15), data_in(15), data_in(15), 
      data_in(15), data_in(15), data_in(15), data_in(14), data_in(13), 
      data_in(12), data_in(11), data_in(10), data_in(9), data_in(8), data_in(7)
      , data_in(6), data_in(5), data_in(4), data_in(3), data_in(2), data_in(1),
      data_in(0) );

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity register_file_nbit_reg32_n_reg32_nbit_addr5 is

   port( reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, add_rd2 
         : in std_logic_vector (4 downto 0);  datain : in std_logic_vector (31 
         downto 0);  out1, out2 : out std_logic_vector (31 downto 0));

end register_file_nbit_reg32_n_reg32_nbit_addr5;

architecture SYN_BEHAVIORAL of register_file_nbit_reg32_n_reg32_nbit_addr5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal registers_1_31_port, registers_1_30_port, registers_1_29_port, 
      registers_1_28_port, registers_1_27_port, registers_1_26_port, 
      registers_1_25_port, registers_1_24_port, registers_1_23_port, 
      registers_1_22_port, registers_1_21_port, registers_1_20_port, 
      registers_1_19_port, registers_1_18_port, registers_1_17_port, 
      registers_1_16_port, registers_1_15_port, registers_1_14_port, 
      registers_1_13_port, registers_1_12_port, registers_1_11_port, 
      registers_1_10_port, registers_1_9_port, registers_1_8_port, 
      registers_1_7_port, registers_1_6_port, registers_1_5_port, 
      registers_1_4_port, registers_1_3_port, registers_1_2_port, 
      registers_1_1_port, registers_1_0_port, registers_2_31_port, 
      registers_2_30_port, registers_2_29_port, registers_2_28_port, 
      registers_2_27_port, registers_2_26_port, registers_2_25_port, 
      registers_2_24_port, registers_2_23_port, registers_2_22_port, 
      registers_2_21_port, registers_2_20_port, registers_2_19_port, 
      registers_2_18_port, registers_2_17_port, registers_2_16_port, 
      registers_2_15_port, registers_2_14_port, registers_2_13_port, 
      registers_2_12_port, registers_2_11_port, registers_2_10_port, 
      registers_2_9_port, registers_2_8_port, registers_2_7_port, 
      registers_2_6_port, registers_2_5_port, registers_2_4_port, 
      registers_2_3_port, registers_2_2_port, registers_2_1_port, 
      registers_2_0_port, registers_3_31_port, registers_3_30_port, 
      registers_3_29_port, registers_3_28_port, registers_3_27_port, 
      registers_3_26_port, registers_3_25_port, registers_3_24_port, 
      registers_3_23_port, registers_3_22_port, registers_3_21_port, 
      registers_3_20_port, registers_3_19_port, registers_3_18_port, 
      registers_3_17_port, registers_3_16_port, registers_3_15_port, 
      registers_3_14_port, registers_3_13_port, registers_3_12_port, 
      registers_3_11_port, registers_3_10_port, registers_3_9_port, 
      registers_3_8_port, registers_3_7_port, registers_3_6_port, 
      registers_3_5_port, registers_3_4_port, registers_3_3_port, 
      registers_3_2_port, registers_3_1_port, registers_3_0_port, 
      registers_4_31_port, registers_4_30_port, registers_4_29_port, 
      registers_4_28_port, registers_4_27_port, registers_4_26_port, 
      registers_4_25_port, registers_4_24_port, registers_4_23_port, 
      registers_4_22_port, registers_4_21_port, registers_4_20_port, 
      registers_4_19_port, registers_4_18_port, registers_4_17_port, 
      registers_4_16_port, registers_4_15_port, registers_4_14_port, 
      registers_4_13_port, registers_4_12_port, registers_4_11_port, 
      registers_4_10_port, registers_4_9_port, registers_4_8_port, 
      registers_4_7_port, registers_4_6_port, registers_4_5_port, 
      registers_4_4_port, registers_4_3_port, registers_4_2_port, 
      registers_4_1_port, registers_4_0_port, registers_5_31_port, 
      registers_5_30_port, registers_5_29_port, registers_5_28_port, 
      registers_5_27_port, registers_5_26_port, registers_5_25_port, 
      registers_5_24_port, registers_5_23_port, registers_5_22_port, 
      registers_5_21_port, registers_5_20_port, registers_5_19_port, 
      registers_5_18_port, registers_5_17_port, registers_5_16_port, 
      registers_5_15_port, registers_5_14_port, registers_5_13_port, 
      registers_5_12_port, registers_5_11_port, registers_5_10_port, 
      registers_5_9_port, registers_5_8_port, registers_5_7_port, 
      registers_5_6_port, registers_5_5_port, registers_5_4_port, 
      registers_5_3_port, registers_5_2_port, registers_5_1_port, 
      registers_5_0_port, registers_6_31_port, registers_6_30_port, 
      registers_6_29_port, registers_6_28_port, registers_6_27_port, 
      registers_6_26_port, registers_6_25_port, registers_6_24_port, 
      registers_6_23_port, registers_6_22_port, registers_6_21_port, 
      registers_6_20_port, registers_6_19_port, registers_6_18_port, 
      registers_6_17_port, registers_6_16_port, registers_6_15_port, 
      registers_6_14_port, registers_6_13_port, registers_6_12_port, 
      registers_6_11_port, registers_6_10_port, registers_6_9_port, 
      registers_6_8_port, registers_6_7_port, registers_6_6_port, 
      registers_6_5_port, registers_6_4_port, registers_6_3_port, 
      registers_6_2_port, registers_6_1_port, registers_6_0_port, 
      registers_7_31_port, registers_7_30_port, registers_7_29_port, 
      registers_7_28_port, registers_7_27_port, registers_7_26_port, 
      registers_7_25_port, registers_7_24_port, registers_7_23_port, 
      registers_7_22_port, registers_7_21_port, registers_7_20_port, 
      registers_7_19_port, registers_7_18_port, registers_7_17_port, 
      registers_7_16_port, registers_7_15_port, registers_7_14_port, 
      registers_7_13_port, registers_7_12_port, registers_7_11_port, 
      registers_7_10_port, registers_7_9_port, registers_7_8_port, 
      registers_7_7_port, registers_7_6_port, registers_7_5_port, 
      registers_7_4_port, registers_7_3_port, registers_7_2_port, 
      registers_7_1_port, registers_7_0_port, registers_8_31_port, 
      registers_8_30_port, registers_8_29_port, registers_8_28_port, 
      registers_8_27_port, registers_8_26_port, registers_8_25_port, 
      registers_8_24_port, registers_8_23_port, registers_8_22_port, 
      registers_8_21_port, registers_8_20_port, registers_8_19_port, 
      registers_8_18_port, registers_8_17_port, registers_8_16_port, 
      registers_8_15_port, registers_8_14_port, registers_8_13_port, 
      registers_8_12_port, registers_8_11_port, registers_8_10_port, 
      registers_8_9_port, registers_8_8_port, registers_8_7_port, 
      registers_8_6_port, registers_8_5_port, registers_8_4_port, 
      registers_8_3_port, registers_8_2_port, registers_8_1_port, 
      registers_8_0_port, registers_9_31_port, registers_9_30_port, 
      registers_9_29_port, registers_9_28_port, registers_9_27_port, 
      registers_9_26_port, registers_9_25_port, registers_9_24_port, 
      registers_9_23_port, registers_9_22_port, registers_9_21_port, 
      registers_9_20_port, registers_9_19_port, registers_9_18_port, 
      registers_9_17_port, registers_9_16_port, registers_9_15_port, 
      registers_9_14_port, registers_9_13_port, registers_9_12_port, 
      registers_9_11_port, registers_9_10_port, registers_9_9_port, 
      registers_9_8_port, registers_9_7_port, registers_9_6_port, 
      registers_9_5_port, registers_9_4_port, registers_9_3_port, 
      registers_9_2_port, registers_9_1_port, registers_9_0_port, 
      registers_10_31_port, registers_10_30_port, registers_10_29_port, 
      registers_10_28_port, registers_10_27_port, registers_10_26_port, 
      registers_10_25_port, registers_10_24_port, registers_10_23_port, 
      registers_10_22_port, registers_10_21_port, registers_10_20_port, 
      registers_10_19_port, registers_10_18_port, registers_10_17_port, 
      registers_10_16_port, registers_10_15_port, registers_10_14_port, 
      registers_10_13_port, registers_10_12_port, registers_10_11_port, 
      registers_10_10_port, registers_10_9_port, registers_10_8_port, 
      registers_10_7_port, registers_10_6_port, registers_10_5_port, 
      registers_10_4_port, registers_10_3_port, registers_10_2_port, 
      registers_10_1_port, registers_10_0_port, registers_11_31_port, 
      registers_11_30_port, registers_11_29_port, registers_11_28_port, 
      registers_11_27_port, registers_11_26_port, registers_11_25_port, 
      registers_11_24_port, registers_11_23_port, registers_11_22_port, 
      registers_11_21_port, registers_11_20_port, registers_11_19_port, 
      registers_11_18_port, registers_11_17_port, registers_11_16_port, 
      registers_11_15_port, registers_11_14_port, registers_11_13_port, 
      registers_11_12_port, registers_11_11_port, registers_11_10_port, 
      registers_11_9_port, registers_11_8_port, registers_11_7_port, 
      registers_11_6_port, registers_11_5_port, registers_11_4_port, 
      registers_11_3_port, registers_11_2_port, registers_11_1_port, 
      registers_11_0_port, registers_12_31_port, registers_12_30_port, 
      registers_12_29_port, registers_12_28_port, registers_12_27_port, 
      registers_12_26_port, registers_12_25_port, registers_12_24_port, 
      registers_12_23_port, registers_12_22_port, registers_12_21_port, 
      registers_12_20_port, registers_12_19_port, registers_12_18_port, 
      registers_12_17_port, registers_12_16_port, registers_12_15_port, 
      registers_12_14_port, registers_12_13_port, registers_12_12_port, 
      registers_12_11_port, registers_12_10_port, registers_12_9_port, 
      registers_12_8_port, registers_12_7_port, registers_12_6_port, 
      registers_12_5_port, registers_12_4_port, registers_12_3_port, 
      registers_12_2_port, registers_12_1_port, registers_12_0_port, 
      registers_13_31_port, registers_13_30_port, registers_13_29_port, 
      registers_13_28_port, registers_13_27_port, registers_13_26_port, 
      registers_13_25_port, registers_13_24_port, registers_13_23_port, 
      registers_13_22_port, registers_13_21_port, registers_13_20_port, 
      registers_13_19_port, registers_13_18_port, registers_13_17_port, 
      registers_13_16_port, registers_13_15_port, registers_13_14_port, 
      registers_13_13_port, registers_13_12_port, registers_13_11_port, 
      registers_13_10_port, registers_13_9_port, registers_13_8_port, 
      registers_13_7_port, registers_13_6_port, registers_13_5_port, 
      registers_13_4_port, registers_13_3_port, registers_13_2_port, 
      registers_13_1_port, registers_13_0_port, registers_14_31_port, 
      registers_14_30_port, registers_14_29_port, registers_14_28_port, 
      registers_14_27_port, registers_14_26_port, registers_14_25_port, 
      registers_14_24_port, registers_14_23_port, registers_14_22_port, 
      registers_14_21_port, registers_14_20_port, registers_14_19_port, 
      registers_14_18_port, registers_14_17_port, registers_14_16_port, 
      registers_14_15_port, registers_14_14_port, registers_14_13_port, 
      registers_14_12_port, registers_14_11_port, registers_14_10_port, 
      registers_14_9_port, registers_14_8_port, registers_14_7_port, 
      registers_14_6_port, registers_14_5_port, registers_14_4_port, 
      registers_14_3_port, registers_14_2_port, registers_14_1_port, 
      registers_14_0_port, registers_15_31_port, registers_15_30_port, 
      registers_15_29_port, registers_15_28_port, registers_15_27_port, 
      registers_15_26_port, registers_15_25_port, registers_15_24_port, 
      registers_15_23_port, registers_15_22_port, registers_15_21_port, 
      registers_15_20_port, registers_15_19_port, registers_15_18_port, 
      registers_15_17_port, registers_15_16_port, registers_15_15_port, 
      registers_15_14_port, registers_15_13_port, registers_15_12_port, 
      registers_15_11_port, registers_15_10_port, registers_15_9_port, 
      registers_15_8_port, registers_15_7_port, registers_15_6_port, 
      registers_15_5_port, registers_15_4_port, registers_15_3_port, 
      registers_15_2_port, registers_15_1_port, registers_15_0_port, 
      registers_16_31_port, registers_16_30_port, registers_16_29_port, 
      registers_16_28_port, registers_16_27_port, registers_16_26_port, 
      registers_16_25_port, registers_16_24_port, registers_16_23_port, 
      registers_16_22_port, registers_16_21_port, registers_16_20_port, 
      registers_16_19_port, registers_16_18_port, registers_16_17_port, 
      registers_16_16_port, registers_16_15_port, registers_16_14_port, 
      registers_16_13_port, registers_16_12_port, registers_16_11_port, 
      registers_16_10_port, registers_16_9_port, registers_16_8_port, 
      registers_16_7_port, registers_16_6_port, registers_16_5_port, 
      registers_16_4_port, registers_16_3_port, registers_16_2_port, 
      registers_16_1_port, registers_16_0_port, registers_17_31_port, 
      registers_17_30_port, registers_17_29_port, registers_17_28_port, 
      registers_17_27_port, registers_17_26_port, registers_17_25_port, 
      registers_17_24_port, registers_17_23_port, registers_17_22_port, 
      registers_17_21_port, registers_17_20_port, registers_17_19_port, 
      registers_17_18_port, registers_17_17_port, registers_17_16_port, 
      registers_17_15_port, registers_17_14_port, registers_17_13_port, 
      registers_17_12_port, registers_17_11_port, registers_17_10_port, 
      registers_17_9_port, registers_17_8_port, registers_17_7_port, 
      registers_17_6_port, registers_17_5_port, registers_17_4_port, 
      registers_17_3_port, registers_17_2_port, registers_17_1_port, 
      registers_17_0_port, registers_18_31_port, registers_18_30_port, 
      registers_18_29_port, registers_18_28_port, registers_18_27_port, 
      registers_18_26_port, registers_18_25_port, registers_18_24_port, 
      registers_18_23_port, registers_18_22_port, registers_18_21_port, 
      registers_18_20_port, registers_18_19_port, registers_18_18_port, 
      registers_18_17_port, registers_18_16_port, registers_18_15_port, 
      registers_18_14_port, registers_18_13_port, registers_18_12_port, 
      registers_18_11_port, registers_18_10_port, registers_18_9_port, 
      registers_18_8_port, registers_18_7_port, registers_18_6_port, 
      registers_18_5_port, registers_18_4_port, registers_18_3_port, 
      registers_18_2_port, registers_18_1_port, registers_18_0_port, 
      registers_19_31_port, registers_19_30_port, registers_19_29_port, 
      registers_19_28_port, registers_19_27_port, registers_19_26_port, 
      registers_19_25_port, registers_19_24_port, registers_19_23_port, 
      registers_19_22_port, registers_19_21_port, registers_19_20_port, 
      registers_19_19_port, registers_19_18_port, registers_19_17_port, 
      registers_19_16_port, registers_19_15_port, registers_19_14_port, 
      registers_19_13_port, registers_19_12_port, registers_19_11_port, 
      registers_19_10_port, registers_19_9_port, registers_19_8_port, 
      registers_19_7_port, registers_19_6_port, registers_19_5_port, 
      registers_19_4_port, registers_19_3_port, registers_19_2_port, 
      registers_19_1_port, registers_19_0_port, registers_20_31_port, 
      registers_20_30_port, registers_20_29_port, registers_20_28_port, 
      registers_20_27_port, registers_20_26_port, registers_20_25_port, 
      registers_20_24_port, registers_20_23_port, registers_20_22_port, 
      registers_20_21_port, registers_20_20_port, registers_20_19_port, 
      registers_20_18_port, registers_20_17_port, registers_20_16_port, 
      registers_20_15_port, registers_20_14_port, registers_20_13_port, 
      registers_20_12_port, registers_20_11_port, registers_20_10_port, 
      registers_20_9_port, registers_20_8_port, registers_20_7_port, 
      registers_20_6_port, registers_20_5_port, registers_20_4_port, 
      registers_20_3_port, registers_20_2_port, registers_20_1_port, 
      registers_20_0_port, registers_21_31_port, registers_21_30_port, 
      registers_21_29_port, registers_21_28_port, registers_21_27_port, 
      registers_21_26_port, registers_21_25_port, registers_21_24_port, 
      registers_21_23_port, registers_21_22_port, registers_21_21_port, 
      registers_21_20_port, registers_21_19_port, registers_21_18_port, 
      registers_21_17_port, registers_21_16_port, registers_21_15_port, 
      registers_21_14_port, registers_21_13_port, registers_21_12_port, 
      registers_21_11_port, registers_21_10_port, registers_21_9_port, 
      registers_21_8_port, registers_21_7_port, registers_21_6_port, 
      registers_21_5_port, registers_21_4_port, registers_21_3_port, 
      registers_21_2_port, registers_21_1_port, registers_21_0_port, 
      registers_22_31_port, registers_22_30_port, registers_22_29_port, 
      registers_22_28_port, registers_22_27_port, registers_22_26_port, 
      registers_22_25_port, registers_22_24_port, registers_22_23_port, 
      registers_22_22_port, registers_22_21_port, registers_22_20_port, 
      registers_22_19_port, registers_22_18_port, registers_22_17_port, 
      registers_22_16_port, registers_22_15_port, registers_22_14_port, 
      registers_22_13_port, registers_22_12_port, registers_22_11_port, 
      registers_22_10_port, registers_22_9_port, registers_22_8_port, 
      registers_22_7_port, registers_22_6_port, registers_22_5_port, 
      registers_22_4_port, registers_22_3_port, registers_22_2_port, 
      registers_22_1_port, registers_22_0_port, registers_23_31_port, 
      registers_23_30_port, registers_23_29_port, registers_23_28_port, 
      registers_23_27_port, registers_23_26_port, registers_23_25_port, 
      registers_23_24_port, registers_23_23_port, registers_23_22_port, 
      registers_23_21_port, registers_23_20_port, registers_23_19_port, 
      registers_23_18_port, registers_23_17_port, registers_23_16_port, 
      registers_23_15_port, registers_23_14_port, registers_23_13_port, 
      registers_23_12_port, registers_23_11_port, registers_23_10_port, 
      registers_23_9_port, registers_23_8_port, registers_23_7_port, 
      registers_23_6_port, registers_23_5_port, registers_23_4_port, 
      registers_23_3_port, registers_23_2_port, registers_23_1_port, 
      registers_23_0_port, registers_24_31_port, registers_24_30_port, 
      registers_24_29_port, registers_24_28_port, registers_24_27_port, 
      registers_24_26_port, registers_24_25_port, registers_24_24_port, 
      registers_24_23_port, registers_24_22_port, registers_24_21_port, 
      registers_24_20_port, registers_24_19_port, registers_24_18_port, 
      registers_24_17_port, registers_24_16_port, registers_24_15_port, 
      registers_24_14_port, registers_24_13_port, registers_24_12_port, 
      registers_24_11_port, registers_24_10_port, registers_24_9_port, 
      registers_24_8_port, registers_24_7_port, registers_24_6_port, 
      registers_24_5_port, registers_24_4_port, registers_24_3_port, 
      registers_24_2_port, registers_24_1_port, registers_24_0_port, 
      registers_25_31_port, registers_25_30_port, registers_25_29_port, 
      registers_25_28_port, registers_25_27_port, registers_25_26_port, 
      registers_25_25_port, registers_25_24_port, registers_25_23_port, 
      registers_25_22_port, registers_25_21_port, registers_25_20_port, 
      registers_25_19_port, registers_25_18_port, registers_25_17_port, 
      registers_25_16_port, registers_25_15_port, registers_25_14_port, 
      registers_25_13_port, registers_25_12_port, registers_25_11_port, 
      registers_25_10_port, registers_25_9_port, registers_25_8_port, 
      registers_25_7_port, registers_25_6_port, registers_25_5_port, 
      registers_25_4_port, registers_25_3_port, registers_25_2_port, 
      registers_25_1_port, registers_25_0_port, registers_26_31_port, 
      registers_26_30_port, registers_26_29_port, registers_26_28_port, 
      registers_26_27_port, registers_26_26_port, registers_26_25_port, 
      registers_26_24_port, registers_26_23_port, registers_26_22_port, 
      registers_26_21_port, registers_26_20_port, registers_26_19_port, 
      registers_26_18_port, registers_26_17_port, registers_26_16_port, 
      registers_26_15_port, registers_26_14_port, registers_26_13_port, 
      registers_26_12_port, registers_26_11_port, registers_26_10_port, 
      registers_26_9_port, registers_26_8_port, registers_26_7_port, 
      registers_26_6_port, registers_26_5_port, registers_26_4_port, 
      registers_26_3_port, registers_26_2_port, registers_26_1_port, 
      registers_26_0_port, registers_27_31_port, registers_27_30_port, 
      registers_27_29_port, registers_27_28_port, registers_27_27_port, 
      registers_27_26_port, registers_27_25_port, registers_27_24_port, 
      registers_27_23_port, registers_27_22_port, registers_27_21_port, 
      registers_27_20_port, registers_27_19_port, registers_27_18_port, 
      registers_27_17_port, registers_27_16_port, registers_27_15_port, 
      registers_27_14_port, registers_27_13_port, registers_27_12_port, 
      registers_27_11_port, registers_27_10_port, registers_27_9_port, 
      registers_27_8_port, registers_27_7_port, registers_27_6_port, 
      registers_27_5_port, registers_27_4_port, registers_27_3_port, 
      registers_27_2_port, registers_27_1_port, registers_27_0_port, 
      registers_28_31_port, registers_28_30_port, registers_28_29_port, 
      registers_28_28_port, registers_28_27_port, registers_28_26_port, 
      registers_28_25_port, registers_28_24_port, registers_28_23_port, 
      registers_28_22_port, registers_28_21_port, registers_28_20_port, 
      registers_28_19_port, registers_28_18_port, registers_28_17_port, 
      registers_28_16_port, registers_28_15_port, registers_28_14_port, 
      registers_28_13_port, registers_28_12_port, registers_28_11_port, 
      registers_28_10_port, registers_28_9_port, registers_28_8_port, 
      registers_28_7_port, registers_28_6_port, registers_28_5_port, 
      registers_28_4_port, registers_28_3_port, registers_28_2_port, 
      registers_28_1_port, registers_28_0_port, registers_29_31_port, 
      registers_29_30_port, registers_29_29_port, registers_29_28_port, 
      registers_29_27_port, registers_29_26_port, registers_29_25_port, 
      registers_29_24_port, registers_29_23_port, registers_29_22_port, 
      registers_29_21_port, registers_29_20_port, registers_29_19_port, 
      registers_29_18_port, registers_29_17_port, registers_29_16_port, 
      registers_29_15_port, registers_29_14_port, registers_29_13_port, 
      registers_29_12_port, registers_29_11_port, registers_29_10_port, 
      registers_29_9_port, registers_29_8_port, registers_29_7_port, 
      registers_29_6_port, registers_29_5_port, registers_29_4_port, 
      registers_29_3_port, registers_29_2_port, registers_29_1_port, 
      registers_29_0_port, registers_30_31_port, registers_30_30_port, 
      registers_30_29_port, registers_30_28_port, registers_30_27_port, 
      registers_30_26_port, registers_30_25_port, registers_30_24_port, 
      registers_30_23_port, registers_30_22_port, registers_30_21_port, 
      registers_30_20_port, registers_30_19_port, registers_30_18_port, 
      registers_30_17_port, registers_30_16_port, registers_30_15_port, 
      registers_30_14_port, registers_30_13_port, registers_30_12_port, 
      registers_30_11_port, registers_30_10_port, registers_30_9_port, 
      registers_30_8_port, registers_30_7_port, registers_30_6_port, 
      registers_30_5_port, registers_30_4_port, registers_30_3_port, 
      registers_30_2_port, registers_30_1_port, registers_30_0_port, 
      registers_31_31_port, registers_31_30_port, registers_31_29_port, 
      registers_31_28_port, registers_31_27_port, registers_31_26_port, 
      registers_31_25_port, registers_31_24_port, registers_31_23_port, 
      registers_31_22_port, registers_31_21_port, registers_31_20_port, 
      registers_31_19_port, registers_31_18_port, registers_31_17_port, 
      registers_31_16_port, registers_31_15_port, registers_31_14_port, 
      registers_31_13_port, registers_31_12_port, registers_31_11_port, 
      registers_31_10_port, registers_31_9_port, registers_31_8_port, 
      registers_31_7_port, registers_31_6_port, registers_31_5_port, 
      registers_31_4_port, registers_31_3_port, registers_31_2_port, 
      registers_31_1_port, registers_31_0_port, N146, N147, N148, N149, N150, 
      N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, 
      N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, 
      N175, N176, N177, N243, N244, N245, N246, N247, N248, N249, N250, N251, 
      N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, 
      N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N307, 
      N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, 
      N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, 
      N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, 
      N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, 
      N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, 
      N368, N369, N371, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, 
      n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, 
      n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, 
      n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, 
      n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
      n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
      n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, 
      n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
      n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, 
      n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
      n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
      n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
      n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
      n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
      n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, 
      n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
      n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
      n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, 
      n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
      n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, 
      n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
      n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, 
      n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
      n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, 
      n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, 
      n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, 
      n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
      n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, 
      n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, 
      n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
      n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
      n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, 
      n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, 
      n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, 
      n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
      n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, 
      n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
      n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, 
      n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, 
      n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, 
      n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, 
      n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
      n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, 
      n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, 
      n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, 
      n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
      n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, 
      n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, 
      n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
      n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
      n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, 
      n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, 
      n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, 
      n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
      n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, 
      n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
      n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, 
      n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, 
      n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, 
      n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
      n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, 
      n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, 
      n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
      n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
      n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
      n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
      n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, 
      n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, 
      n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, 
      n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, 
      n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, 
      n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, 
      n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, 
      n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
      n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, 
      n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
      n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, 
      n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, 
      n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, 
      n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
      n2685, n2686, n2687, n2688, n2689 : std_logic;

begin
   
   registers_reg_1_31_inst : DLH_X1 port map( G => n1970, D => n2060, Q => 
                           registers_1_31_port);
   registers_reg_1_30_inst : DLH_X1 port map( G => n1970, D => n2063, Q => 
                           registers_1_30_port);
   registers_reg_1_29_inst : DLH_X1 port map( G => n1970, D => n2066, Q => 
                           registers_1_29_port);
   registers_reg_1_28_inst : DLH_X1 port map( G => n1970, D => n2069, Q => 
                           registers_1_28_port);
   registers_reg_1_27_inst : DLH_X1 port map( G => n1970, D => n2072, Q => 
                           registers_1_27_port);
   registers_reg_1_26_inst : DLH_X1 port map( G => n1970, D => n2075, Q => 
                           registers_1_26_port);
   registers_reg_1_25_inst : DLH_X1 port map( G => n1970, D => n2078, Q => 
                           registers_1_25_port);
   registers_reg_1_24_inst : DLH_X1 port map( G => n1969, D => n2081, Q => 
                           registers_1_24_port);
   registers_reg_1_23_inst : DLH_X1 port map( G => n1969, D => n2084, Q => 
                           registers_1_23_port);
   registers_reg_1_22_inst : DLH_X1 port map( G => n1969, D => n2087, Q => 
                           registers_1_22_port);
   registers_reg_1_21_inst : DLH_X1 port map( G => n1969, D => n2090, Q => 
                           registers_1_21_port);
   registers_reg_1_20_inst : DLH_X1 port map( G => n1970, D => n2093, Q => 
                           registers_1_20_port);
   registers_reg_1_19_inst : DLH_X1 port map( G => n1969, D => n2096, Q => 
                           registers_1_19_port);
   registers_reg_1_18_inst : DLH_X1 port map( G => n1969, D => n2099, Q => 
                           registers_1_18_port);
   registers_reg_1_17_inst : DLH_X1 port map( G => n1970, D => n2102, Q => 
                           registers_1_17_port);
   registers_reg_1_16_inst : DLH_X1 port map( G => n1969, D => n2105, Q => 
                           registers_1_16_port);
   registers_reg_1_15_inst : DLH_X1 port map( G => n1969, D => n2108, Q => 
                           registers_1_15_port);
   registers_reg_1_14_inst : DLH_X1 port map( G => n1969, D => n2111, Q => 
                           registers_1_14_port);
   registers_reg_1_13_inst : DLH_X1 port map( G => n1968, D => n2114, Q => 
                           registers_1_13_port);
   registers_reg_1_12_inst : DLH_X1 port map( G => n1969, D => n2117, Q => 
                           registers_1_12_port);
   registers_reg_1_11_inst : DLH_X1 port map( G => n1968, D => n2120, Q => 
                           registers_1_11_port);
   registers_reg_1_10_inst : DLH_X1 port map( G => n1968, D => n2123, Q => 
                           registers_1_10_port);
   registers_reg_1_9_inst : DLH_X1 port map( G => n1968, D => n2126, Q => 
                           registers_1_9_port);
   registers_reg_1_8_inst : DLH_X1 port map( G => n1968, D => n2129, Q => 
                           registers_1_8_port);
   registers_reg_1_7_inst : DLH_X1 port map( G => n1968, D => n2132, Q => 
                           registers_1_7_port);
   registers_reg_1_6_inst : DLH_X1 port map( G => n1968, D => n2135, Q => 
                           registers_1_6_port);
   registers_reg_1_5_inst : DLH_X1 port map( G => n1968, D => n2138, Q => 
                           registers_1_5_port);
   registers_reg_1_4_inst : DLH_X1 port map( G => n1968, D => n2141, Q => 
                           registers_1_4_port);
   registers_reg_1_3_inst : DLH_X1 port map( G => n1968, D => n2144, Q => 
                           registers_1_3_port);
   registers_reg_1_2_inst : DLH_X1 port map( G => n1968, D => n2147, Q => 
                           registers_1_2_port);
   registers_reg_1_1_inst : DLH_X1 port map( G => n1969, D => n2150, Q => 
                           registers_1_1_port);
   registers_reg_1_0_inst : DLH_X1 port map( G => n1970, D => n2153, Q => 
                           registers_1_0_port);
   registers_reg_2_31_inst : DLH_X1 port map( G => n1973, D => n2060, Q => 
                           registers_2_31_port);
   registers_reg_2_30_inst : DLH_X1 port map( G => n1973, D => n2063, Q => 
                           registers_2_30_port);
   registers_reg_2_29_inst : DLH_X1 port map( G => n1973, D => n2066, Q => 
                           registers_2_29_port);
   registers_reg_2_28_inst : DLH_X1 port map( G => n1973, D => n2069, Q => 
                           registers_2_28_port);
   registers_reg_2_27_inst : DLH_X1 port map( G => n1973, D => n2072, Q => 
                           registers_2_27_port);
   registers_reg_2_26_inst : DLH_X1 port map( G => n1973, D => n2075, Q => 
                           registers_2_26_port);
   registers_reg_2_25_inst : DLH_X1 port map( G => n1973, D => n2078, Q => 
                           registers_2_25_port);
   registers_reg_2_24_inst : DLH_X1 port map( G => n1972, D => n2081, Q => 
                           registers_2_24_port);
   registers_reg_2_23_inst : DLH_X1 port map( G => n1972, D => n2084, Q => 
                           registers_2_23_port);
   registers_reg_2_22_inst : DLH_X1 port map( G => n1972, D => n2087, Q => 
                           registers_2_22_port);
   registers_reg_2_21_inst : DLH_X1 port map( G => n1972, D => n2090, Q => 
                           registers_2_21_port);
   registers_reg_2_20_inst : DLH_X1 port map( G => n1973, D => n2093, Q => 
                           registers_2_20_port);
   registers_reg_2_19_inst : DLH_X1 port map( G => n1972, D => n2096, Q => 
                           registers_2_19_port);
   registers_reg_2_18_inst : DLH_X1 port map( G => n1972, D => n2099, Q => 
                           registers_2_18_port);
   registers_reg_2_17_inst : DLH_X1 port map( G => n1973, D => n2102, Q => 
                           registers_2_17_port);
   registers_reg_2_16_inst : DLH_X1 port map( G => n1972, D => n2105, Q => 
                           registers_2_16_port);
   registers_reg_2_15_inst : DLH_X1 port map( G => n1972, D => n2108, Q => 
                           registers_2_15_port);
   registers_reg_2_14_inst : DLH_X1 port map( G => n1972, D => n2111, Q => 
                           registers_2_14_port);
   registers_reg_2_13_inst : DLH_X1 port map( G => n1971, D => n2114, Q => 
                           registers_2_13_port);
   registers_reg_2_12_inst : DLH_X1 port map( G => n1972, D => n2117, Q => 
                           registers_2_12_port);
   registers_reg_2_11_inst : DLH_X1 port map( G => n1971, D => n2120, Q => 
                           registers_2_11_port);
   registers_reg_2_10_inst : DLH_X1 port map( G => n1971, D => n2123, Q => 
                           registers_2_10_port);
   registers_reg_2_9_inst : DLH_X1 port map( G => n1971, D => n2126, Q => 
                           registers_2_9_port);
   registers_reg_2_8_inst : DLH_X1 port map( G => n1971, D => n2129, Q => 
                           registers_2_8_port);
   registers_reg_2_7_inst : DLH_X1 port map( G => n1971, D => n2132, Q => 
                           registers_2_7_port);
   registers_reg_2_6_inst : DLH_X1 port map( G => n1971, D => n2135, Q => 
                           registers_2_6_port);
   registers_reg_2_5_inst : DLH_X1 port map( G => n1971, D => n2138, Q => 
                           registers_2_5_port);
   registers_reg_2_4_inst : DLH_X1 port map( G => n1971, D => n2141, Q => 
                           registers_2_4_port);
   registers_reg_2_3_inst : DLH_X1 port map( G => n1971, D => n2144, Q => 
                           registers_2_3_port);
   registers_reg_2_2_inst : DLH_X1 port map( G => n1971, D => n2147, Q => 
                           registers_2_2_port);
   registers_reg_2_1_inst : DLH_X1 port map( G => n1972, D => n2150, Q => 
                           registers_2_1_port);
   registers_reg_2_0_inst : DLH_X1 port map( G => n1973, D => n2153, Q => 
                           registers_2_0_port);
   registers_reg_3_31_inst : DLH_X1 port map( G => n1976, D => n2060, Q => 
                           registers_3_31_port);
   registers_reg_3_30_inst : DLH_X1 port map( G => n1976, D => n2063, Q => 
                           registers_3_30_port);
   registers_reg_3_29_inst : DLH_X1 port map( G => n1976, D => n2066, Q => 
                           registers_3_29_port);
   registers_reg_3_28_inst : DLH_X1 port map( G => n1976, D => n2069, Q => 
                           registers_3_28_port);
   registers_reg_3_27_inst : DLH_X1 port map( G => n1976, D => n2072, Q => 
                           registers_3_27_port);
   registers_reg_3_26_inst : DLH_X1 port map( G => n1976, D => n2075, Q => 
                           registers_3_26_port);
   registers_reg_3_25_inst : DLH_X1 port map( G => n1976, D => n2078, Q => 
                           registers_3_25_port);
   registers_reg_3_24_inst : DLH_X1 port map( G => n1975, D => n2081, Q => 
                           registers_3_24_port);
   registers_reg_3_23_inst : DLH_X1 port map( G => n1975, D => n2084, Q => 
                           registers_3_23_port);
   registers_reg_3_22_inst : DLH_X1 port map( G => n1975, D => n2087, Q => 
                           registers_3_22_port);
   registers_reg_3_21_inst : DLH_X1 port map( G => n1975, D => n2090, Q => 
                           registers_3_21_port);
   registers_reg_3_20_inst : DLH_X1 port map( G => n1976, D => n2093, Q => 
                           registers_3_20_port);
   registers_reg_3_19_inst : DLH_X1 port map( G => n1975, D => n2096, Q => 
                           registers_3_19_port);
   registers_reg_3_18_inst : DLH_X1 port map( G => n1975, D => n2099, Q => 
                           registers_3_18_port);
   registers_reg_3_17_inst : DLH_X1 port map( G => n1976, D => n2102, Q => 
                           registers_3_17_port);
   registers_reg_3_16_inst : DLH_X1 port map( G => n1975, D => n2105, Q => 
                           registers_3_16_port);
   registers_reg_3_15_inst : DLH_X1 port map( G => n1975, D => n2108, Q => 
                           registers_3_15_port);
   registers_reg_3_14_inst : DLH_X1 port map( G => n1975, D => n2111, Q => 
                           registers_3_14_port);
   registers_reg_3_13_inst : DLH_X1 port map( G => n1974, D => n2114, Q => 
                           registers_3_13_port);
   registers_reg_3_12_inst : DLH_X1 port map( G => n1975, D => n2117, Q => 
                           registers_3_12_port);
   registers_reg_3_11_inst : DLH_X1 port map( G => n1974, D => n2120, Q => 
                           registers_3_11_port);
   registers_reg_3_10_inst : DLH_X1 port map( G => n1974, D => n2123, Q => 
                           registers_3_10_port);
   registers_reg_3_9_inst : DLH_X1 port map( G => n1974, D => n2126, Q => 
                           registers_3_9_port);
   registers_reg_3_8_inst : DLH_X1 port map( G => n1974, D => n2129, Q => 
                           registers_3_8_port);
   registers_reg_3_7_inst : DLH_X1 port map( G => n1974, D => n2132, Q => 
                           registers_3_7_port);
   registers_reg_3_6_inst : DLH_X1 port map( G => n1974, D => n2135, Q => 
                           registers_3_6_port);
   registers_reg_3_5_inst : DLH_X1 port map( G => n1974, D => n2138, Q => 
                           registers_3_5_port);
   registers_reg_3_4_inst : DLH_X1 port map( G => n1974, D => n2141, Q => 
                           registers_3_4_port);
   registers_reg_3_3_inst : DLH_X1 port map( G => n1974, D => n2144, Q => 
                           registers_3_3_port);
   registers_reg_3_2_inst : DLH_X1 port map( G => n1974, D => n2147, Q => 
                           registers_3_2_port);
   registers_reg_3_1_inst : DLH_X1 port map( G => n1975, D => n2150, Q => 
                           registers_3_1_port);
   registers_reg_3_0_inst : DLH_X1 port map( G => n1976, D => n2153, Q => 
                           registers_3_0_port);
   registers_reg_4_31_inst : DLH_X1 port map( G => n1979, D => n2060, Q => 
                           registers_4_31_port);
   registers_reg_4_30_inst : DLH_X1 port map( G => n1979, D => n2063, Q => 
                           registers_4_30_port);
   registers_reg_4_29_inst : DLH_X1 port map( G => n1979, D => n2066, Q => 
                           registers_4_29_port);
   registers_reg_4_28_inst : DLH_X1 port map( G => n1979, D => n2069, Q => 
                           registers_4_28_port);
   registers_reg_4_27_inst : DLH_X1 port map( G => n1979, D => n2072, Q => 
                           registers_4_27_port);
   registers_reg_4_26_inst : DLH_X1 port map( G => n1979, D => n2075, Q => 
                           registers_4_26_port);
   registers_reg_4_25_inst : DLH_X1 port map( G => n1979, D => n2078, Q => 
                           registers_4_25_port);
   registers_reg_4_24_inst : DLH_X1 port map( G => n1978, D => n2081, Q => 
                           registers_4_24_port);
   registers_reg_4_23_inst : DLH_X1 port map( G => n1978, D => n2084, Q => 
                           registers_4_23_port);
   registers_reg_4_22_inst : DLH_X1 port map( G => n1978, D => n2087, Q => 
                           registers_4_22_port);
   registers_reg_4_21_inst : DLH_X1 port map( G => n1978, D => n2090, Q => 
                           registers_4_21_port);
   registers_reg_4_20_inst : DLH_X1 port map( G => n1979, D => n2093, Q => 
                           registers_4_20_port);
   registers_reg_4_19_inst : DLH_X1 port map( G => n1978, D => n2096, Q => 
                           registers_4_19_port);
   registers_reg_4_18_inst : DLH_X1 port map( G => n1978, D => n2099, Q => 
                           registers_4_18_port);
   registers_reg_4_17_inst : DLH_X1 port map( G => n1979, D => n2102, Q => 
                           registers_4_17_port);
   registers_reg_4_16_inst : DLH_X1 port map( G => n1978, D => n2105, Q => 
                           registers_4_16_port);
   registers_reg_4_15_inst : DLH_X1 port map( G => n1978, D => n2108, Q => 
                           registers_4_15_port);
   registers_reg_4_14_inst : DLH_X1 port map( G => n1978, D => n2111, Q => 
                           registers_4_14_port);
   registers_reg_4_13_inst : DLH_X1 port map( G => n1977, D => n2114, Q => 
                           registers_4_13_port);
   registers_reg_4_12_inst : DLH_X1 port map( G => n1978, D => n2117, Q => 
                           registers_4_12_port);
   registers_reg_4_11_inst : DLH_X1 port map( G => n1977, D => n2120, Q => 
                           registers_4_11_port);
   registers_reg_4_10_inst : DLH_X1 port map( G => n1977, D => n2123, Q => 
                           registers_4_10_port);
   registers_reg_4_9_inst : DLH_X1 port map( G => n1977, D => n2126, Q => 
                           registers_4_9_port);
   registers_reg_4_8_inst : DLH_X1 port map( G => n1977, D => n2129, Q => 
                           registers_4_8_port);
   registers_reg_4_7_inst : DLH_X1 port map( G => n1977, D => n2132, Q => 
                           registers_4_7_port);
   registers_reg_4_6_inst : DLH_X1 port map( G => n1977, D => n2135, Q => 
                           registers_4_6_port);
   registers_reg_4_5_inst : DLH_X1 port map( G => n1977, D => n2138, Q => 
                           registers_4_5_port);
   registers_reg_4_4_inst : DLH_X1 port map( G => n1977, D => n2141, Q => 
                           registers_4_4_port);
   registers_reg_4_3_inst : DLH_X1 port map( G => n1977, D => n2144, Q => 
                           registers_4_3_port);
   registers_reg_4_2_inst : DLH_X1 port map( G => n1977, D => n2147, Q => 
                           registers_4_2_port);
   registers_reg_4_1_inst : DLH_X1 port map( G => n1978, D => n2150, Q => 
                           registers_4_1_port);
   registers_reg_4_0_inst : DLH_X1 port map( G => n1979, D => n2153, Q => 
                           registers_4_0_port);
   registers_reg_5_31_inst : DLH_X1 port map( G => n1982, D => n2060, Q => 
                           registers_5_31_port);
   registers_reg_5_30_inst : DLH_X1 port map( G => n1982, D => n2063, Q => 
                           registers_5_30_port);
   registers_reg_5_29_inst : DLH_X1 port map( G => n1982, D => n2066, Q => 
                           registers_5_29_port);
   registers_reg_5_28_inst : DLH_X1 port map( G => n1982, D => n2069, Q => 
                           registers_5_28_port);
   registers_reg_5_27_inst : DLH_X1 port map( G => n1982, D => n2072, Q => 
                           registers_5_27_port);
   registers_reg_5_26_inst : DLH_X1 port map( G => n1982, D => n2075, Q => 
                           registers_5_26_port);
   registers_reg_5_25_inst : DLH_X1 port map( G => n1982, D => n2078, Q => 
                           registers_5_25_port);
   registers_reg_5_24_inst : DLH_X1 port map( G => n1981, D => n2081, Q => 
                           registers_5_24_port);
   registers_reg_5_23_inst : DLH_X1 port map( G => n1981, D => n2084, Q => 
                           registers_5_23_port);
   registers_reg_5_22_inst : DLH_X1 port map( G => n1981, D => n2087, Q => 
                           registers_5_22_port);
   registers_reg_5_21_inst : DLH_X1 port map( G => n1981, D => n2090, Q => 
                           registers_5_21_port);
   registers_reg_5_20_inst : DLH_X1 port map( G => n1982, D => n2093, Q => 
                           registers_5_20_port);
   registers_reg_5_19_inst : DLH_X1 port map( G => n1981, D => n2096, Q => 
                           registers_5_19_port);
   registers_reg_5_18_inst : DLH_X1 port map( G => n1981, D => n2099, Q => 
                           registers_5_18_port);
   registers_reg_5_17_inst : DLH_X1 port map( G => n1982, D => n2102, Q => 
                           registers_5_17_port);
   registers_reg_5_16_inst : DLH_X1 port map( G => n1981, D => n2105, Q => 
                           registers_5_16_port);
   registers_reg_5_15_inst : DLH_X1 port map( G => n1981, D => n2108, Q => 
                           registers_5_15_port);
   registers_reg_5_14_inst : DLH_X1 port map( G => n1981, D => n2111, Q => 
                           registers_5_14_port);
   registers_reg_5_13_inst : DLH_X1 port map( G => n1980, D => n2114, Q => 
                           registers_5_13_port);
   registers_reg_5_12_inst : DLH_X1 port map( G => n1981, D => n2117, Q => 
                           registers_5_12_port);
   registers_reg_5_11_inst : DLH_X1 port map( G => n1980, D => n2120, Q => 
                           registers_5_11_port);
   registers_reg_5_10_inst : DLH_X1 port map( G => n1980, D => n2123, Q => 
                           registers_5_10_port);
   registers_reg_5_9_inst : DLH_X1 port map( G => n1980, D => n2126, Q => 
                           registers_5_9_port);
   registers_reg_5_8_inst : DLH_X1 port map( G => n1980, D => n2129, Q => 
                           registers_5_8_port);
   registers_reg_5_7_inst : DLH_X1 port map( G => n1980, D => n2132, Q => 
                           registers_5_7_port);
   registers_reg_5_6_inst : DLH_X1 port map( G => n1980, D => n2135, Q => 
                           registers_5_6_port);
   registers_reg_5_5_inst : DLH_X1 port map( G => n1980, D => n2138, Q => 
                           registers_5_5_port);
   registers_reg_5_4_inst : DLH_X1 port map( G => n1980, D => n2141, Q => 
                           registers_5_4_port);
   registers_reg_5_3_inst : DLH_X1 port map( G => n1980, D => n2144, Q => 
                           registers_5_3_port);
   registers_reg_5_2_inst : DLH_X1 port map( G => n1980, D => n2147, Q => 
                           registers_5_2_port);
   registers_reg_5_1_inst : DLH_X1 port map( G => n1981, D => n2150, Q => 
                           registers_5_1_port);
   registers_reg_5_0_inst : DLH_X1 port map( G => n1982, D => n2153, Q => 
                           registers_5_0_port);
   registers_reg_6_31_inst : DLH_X1 port map( G => n1985, D => n2060, Q => 
                           registers_6_31_port);
   registers_reg_6_30_inst : DLH_X1 port map( G => n1985, D => n2063, Q => 
                           registers_6_30_port);
   registers_reg_6_29_inst : DLH_X1 port map( G => n1985, D => n2066, Q => 
                           registers_6_29_port);
   registers_reg_6_28_inst : DLH_X1 port map( G => n1985, D => n2069, Q => 
                           registers_6_28_port);
   registers_reg_6_27_inst : DLH_X1 port map( G => n1985, D => n2072, Q => 
                           registers_6_27_port);
   registers_reg_6_26_inst : DLH_X1 port map( G => n1985, D => n2075, Q => 
                           registers_6_26_port);
   registers_reg_6_25_inst : DLH_X1 port map( G => n1985, D => n2078, Q => 
                           registers_6_25_port);
   registers_reg_6_24_inst : DLH_X1 port map( G => n1984, D => n2081, Q => 
                           registers_6_24_port);
   registers_reg_6_23_inst : DLH_X1 port map( G => n1984, D => n2084, Q => 
                           registers_6_23_port);
   registers_reg_6_22_inst : DLH_X1 port map( G => n1984, D => n2087, Q => 
                           registers_6_22_port);
   registers_reg_6_21_inst : DLH_X1 port map( G => n1984, D => n2090, Q => 
                           registers_6_21_port);
   registers_reg_6_20_inst : DLH_X1 port map( G => n1985, D => n2093, Q => 
                           registers_6_20_port);
   registers_reg_6_19_inst : DLH_X1 port map( G => n1984, D => n2096, Q => 
                           registers_6_19_port);
   registers_reg_6_18_inst : DLH_X1 port map( G => n1984, D => n2099, Q => 
                           registers_6_18_port);
   registers_reg_6_17_inst : DLH_X1 port map( G => n1985, D => n2102, Q => 
                           registers_6_17_port);
   registers_reg_6_16_inst : DLH_X1 port map( G => n1984, D => n2105, Q => 
                           registers_6_16_port);
   registers_reg_6_15_inst : DLH_X1 port map( G => n1984, D => n2108, Q => 
                           registers_6_15_port);
   registers_reg_6_14_inst : DLH_X1 port map( G => n1984, D => n2111, Q => 
                           registers_6_14_port);
   registers_reg_6_13_inst : DLH_X1 port map( G => n1983, D => n2114, Q => 
                           registers_6_13_port);
   registers_reg_6_12_inst : DLH_X1 port map( G => n1984, D => n2117, Q => 
                           registers_6_12_port);
   registers_reg_6_11_inst : DLH_X1 port map( G => n1983, D => n2120, Q => 
                           registers_6_11_port);
   registers_reg_6_10_inst : DLH_X1 port map( G => n1983, D => n2123, Q => 
                           registers_6_10_port);
   registers_reg_6_9_inst : DLH_X1 port map( G => n1983, D => n2126, Q => 
                           registers_6_9_port);
   registers_reg_6_8_inst : DLH_X1 port map( G => n1983, D => n2129, Q => 
                           registers_6_8_port);
   registers_reg_6_7_inst : DLH_X1 port map( G => n1983, D => n2132, Q => 
                           registers_6_7_port);
   registers_reg_6_6_inst : DLH_X1 port map( G => n1983, D => n2135, Q => 
                           registers_6_6_port);
   registers_reg_6_5_inst : DLH_X1 port map( G => n1983, D => n2138, Q => 
                           registers_6_5_port);
   registers_reg_6_4_inst : DLH_X1 port map( G => n1983, D => n2141, Q => 
                           registers_6_4_port);
   registers_reg_6_3_inst : DLH_X1 port map( G => n1983, D => n2144, Q => 
                           registers_6_3_port);
   registers_reg_6_2_inst : DLH_X1 port map( G => n1983, D => n2147, Q => 
                           registers_6_2_port);
   registers_reg_6_1_inst : DLH_X1 port map( G => n1984, D => n2150, Q => 
                           registers_6_1_port);
   registers_reg_6_0_inst : DLH_X1 port map( G => n1985, D => n2153, Q => 
                           registers_6_0_port);
   registers_reg_7_31_inst : DLH_X1 port map( G => n1988, D => n2060, Q => 
                           registers_7_31_port);
   registers_reg_7_30_inst : DLH_X1 port map( G => n1988, D => n2063, Q => 
                           registers_7_30_port);
   registers_reg_7_29_inst : DLH_X1 port map( G => n1988, D => n2066, Q => 
                           registers_7_29_port);
   registers_reg_7_28_inst : DLH_X1 port map( G => n1988, D => n2069, Q => 
                           registers_7_28_port);
   registers_reg_7_27_inst : DLH_X1 port map( G => n1988, D => n2072, Q => 
                           registers_7_27_port);
   registers_reg_7_26_inst : DLH_X1 port map( G => n1988, D => n2075, Q => 
                           registers_7_26_port);
   registers_reg_7_25_inst : DLH_X1 port map( G => n1988, D => n2078, Q => 
                           registers_7_25_port);
   registers_reg_7_24_inst : DLH_X1 port map( G => n1987, D => n2081, Q => 
                           registers_7_24_port);
   registers_reg_7_23_inst : DLH_X1 port map( G => n1987, D => n2084, Q => 
                           registers_7_23_port);
   registers_reg_7_22_inst : DLH_X1 port map( G => n1987, D => n2087, Q => 
                           registers_7_22_port);
   registers_reg_7_21_inst : DLH_X1 port map( G => n1987, D => n2090, Q => 
                           registers_7_21_port);
   registers_reg_7_20_inst : DLH_X1 port map( G => n1988, D => n2093, Q => 
                           registers_7_20_port);
   registers_reg_7_19_inst : DLH_X1 port map( G => n1987, D => n2096, Q => 
                           registers_7_19_port);
   registers_reg_7_18_inst : DLH_X1 port map( G => n1987, D => n2099, Q => 
                           registers_7_18_port);
   registers_reg_7_17_inst : DLH_X1 port map( G => n1988, D => n2102, Q => 
                           registers_7_17_port);
   registers_reg_7_16_inst : DLH_X1 port map( G => n1987, D => n2105, Q => 
                           registers_7_16_port);
   registers_reg_7_15_inst : DLH_X1 port map( G => n1987, D => n2108, Q => 
                           registers_7_15_port);
   registers_reg_7_14_inst : DLH_X1 port map( G => n1987, D => n2111, Q => 
                           registers_7_14_port);
   registers_reg_7_13_inst : DLH_X1 port map( G => n1986, D => n2114, Q => 
                           registers_7_13_port);
   registers_reg_7_12_inst : DLH_X1 port map( G => n1987, D => n2117, Q => 
                           registers_7_12_port);
   registers_reg_7_11_inst : DLH_X1 port map( G => n1986, D => n2120, Q => 
                           registers_7_11_port);
   registers_reg_7_10_inst : DLH_X1 port map( G => n1986, D => n2123, Q => 
                           registers_7_10_port);
   registers_reg_7_9_inst : DLH_X1 port map( G => n1986, D => n2126, Q => 
                           registers_7_9_port);
   registers_reg_7_8_inst : DLH_X1 port map( G => n1986, D => n2129, Q => 
                           registers_7_8_port);
   registers_reg_7_7_inst : DLH_X1 port map( G => n1986, D => n2132, Q => 
                           registers_7_7_port);
   registers_reg_7_6_inst : DLH_X1 port map( G => n1986, D => n2135, Q => 
                           registers_7_6_port);
   registers_reg_7_5_inst : DLH_X1 port map( G => n1986, D => n2138, Q => 
                           registers_7_5_port);
   registers_reg_7_4_inst : DLH_X1 port map( G => n1986, D => n2141, Q => 
                           registers_7_4_port);
   registers_reg_7_3_inst : DLH_X1 port map( G => n1986, D => n2144, Q => 
                           registers_7_3_port);
   registers_reg_7_2_inst : DLH_X1 port map( G => n1986, D => n2147, Q => 
                           registers_7_2_port);
   registers_reg_7_1_inst : DLH_X1 port map( G => n1987, D => n2150, Q => 
                           registers_7_1_port);
   registers_reg_7_0_inst : DLH_X1 port map( G => n1988, D => n2153, Q => 
                           registers_7_0_port);
   registers_reg_8_31_inst : DLH_X1 port map( G => n1991, D => n2060, Q => 
                           registers_8_31_port);
   registers_reg_8_30_inst : DLH_X1 port map( G => n1991, D => n2063, Q => 
                           registers_8_30_port);
   registers_reg_8_29_inst : DLH_X1 port map( G => n1991, D => n2066, Q => 
                           registers_8_29_port);
   registers_reg_8_28_inst : DLH_X1 port map( G => n1991, D => n2069, Q => 
                           registers_8_28_port);
   registers_reg_8_27_inst : DLH_X1 port map( G => n1991, D => n2072, Q => 
                           registers_8_27_port);
   registers_reg_8_26_inst : DLH_X1 port map( G => n1991, D => n2075, Q => 
                           registers_8_26_port);
   registers_reg_8_25_inst : DLH_X1 port map( G => n1991, D => n2078, Q => 
                           registers_8_25_port);
   registers_reg_8_24_inst : DLH_X1 port map( G => n1990, D => n2081, Q => 
                           registers_8_24_port);
   registers_reg_8_23_inst : DLH_X1 port map( G => n1990, D => n2084, Q => 
                           registers_8_23_port);
   registers_reg_8_22_inst : DLH_X1 port map( G => n1990, D => n2087, Q => 
                           registers_8_22_port);
   registers_reg_8_21_inst : DLH_X1 port map( G => n1990, D => n2090, Q => 
                           registers_8_21_port);
   registers_reg_8_20_inst : DLH_X1 port map( G => n1991, D => n2093, Q => 
                           registers_8_20_port);
   registers_reg_8_19_inst : DLH_X1 port map( G => n1990, D => n2096, Q => 
                           registers_8_19_port);
   registers_reg_8_18_inst : DLH_X1 port map( G => n1990, D => n2099, Q => 
                           registers_8_18_port);
   registers_reg_8_17_inst : DLH_X1 port map( G => n1991, D => n2102, Q => 
                           registers_8_17_port);
   registers_reg_8_16_inst : DLH_X1 port map( G => n1990, D => n2105, Q => 
                           registers_8_16_port);
   registers_reg_8_15_inst : DLH_X1 port map( G => n1990, D => n2108, Q => 
                           registers_8_15_port);
   registers_reg_8_14_inst : DLH_X1 port map( G => n1990, D => n2111, Q => 
                           registers_8_14_port);
   registers_reg_8_13_inst : DLH_X1 port map( G => n1989, D => n2114, Q => 
                           registers_8_13_port);
   registers_reg_8_12_inst : DLH_X1 port map( G => n1990, D => n2117, Q => 
                           registers_8_12_port);
   registers_reg_8_11_inst : DLH_X1 port map( G => n1989, D => n2120, Q => 
                           registers_8_11_port);
   registers_reg_8_10_inst : DLH_X1 port map( G => n1989, D => n2123, Q => 
                           registers_8_10_port);
   registers_reg_8_9_inst : DLH_X1 port map( G => n1989, D => n2126, Q => 
                           registers_8_9_port);
   registers_reg_8_8_inst : DLH_X1 port map( G => n1989, D => n2129, Q => 
                           registers_8_8_port);
   registers_reg_8_7_inst : DLH_X1 port map( G => n1989, D => n2132, Q => 
                           registers_8_7_port);
   registers_reg_8_6_inst : DLH_X1 port map( G => n1989, D => n2135, Q => 
                           registers_8_6_port);
   registers_reg_8_5_inst : DLH_X1 port map( G => n1989, D => n2138, Q => 
                           registers_8_5_port);
   registers_reg_8_4_inst : DLH_X1 port map( G => n1989, D => n2141, Q => 
                           registers_8_4_port);
   registers_reg_8_3_inst : DLH_X1 port map( G => n1989, D => n2144, Q => 
                           registers_8_3_port);
   registers_reg_8_2_inst : DLH_X1 port map( G => n1989, D => n2147, Q => 
                           registers_8_2_port);
   registers_reg_8_1_inst : DLH_X1 port map( G => n1990, D => n2150, Q => 
                           registers_8_1_port);
   registers_reg_8_0_inst : DLH_X1 port map( G => n1991, D => n2153, Q => 
                           registers_8_0_port);
   registers_reg_9_31_inst : DLH_X1 port map( G => n1994, D => n2060, Q => 
                           registers_9_31_port);
   registers_reg_9_30_inst : DLH_X1 port map( G => n1994, D => n2063, Q => 
                           registers_9_30_port);
   registers_reg_9_29_inst : DLH_X1 port map( G => n1994, D => n2066, Q => 
                           registers_9_29_port);
   registers_reg_9_28_inst : DLH_X1 port map( G => n1994, D => n2069, Q => 
                           registers_9_28_port);
   registers_reg_9_27_inst : DLH_X1 port map( G => n1994, D => n2072, Q => 
                           registers_9_27_port);
   registers_reg_9_26_inst : DLH_X1 port map( G => n1994, D => n2075, Q => 
                           registers_9_26_port);
   registers_reg_9_25_inst : DLH_X1 port map( G => n1994, D => n2078, Q => 
                           registers_9_25_port);
   registers_reg_9_24_inst : DLH_X1 port map( G => n1993, D => n2081, Q => 
                           registers_9_24_port);
   registers_reg_9_23_inst : DLH_X1 port map( G => n1993, D => n2084, Q => 
                           registers_9_23_port);
   registers_reg_9_22_inst : DLH_X1 port map( G => n1993, D => n2087, Q => 
                           registers_9_22_port);
   registers_reg_9_21_inst : DLH_X1 port map( G => n1993, D => n2090, Q => 
                           registers_9_21_port);
   registers_reg_9_20_inst : DLH_X1 port map( G => n1994, D => n2093, Q => 
                           registers_9_20_port);
   registers_reg_9_19_inst : DLH_X1 port map( G => n1993, D => n2096, Q => 
                           registers_9_19_port);
   registers_reg_9_18_inst : DLH_X1 port map( G => n1993, D => n2099, Q => 
                           registers_9_18_port);
   registers_reg_9_17_inst : DLH_X1 port map( G => n1994, D => n2102, Q => 
                           registers_9_17_port);
   registers_reg_9_16_inst : DLH_X1 port map( G => n1993, D => n2105, Q => 
                           registers_9_16_port);
   registers_reg_9_15_inst : DLH_X1 port map( G => n1993, D => n2108, Q => 
                           registers_9_15_port);
   registers_reg_9_14_inst : DLH_X1 port map( G => n1993, D => n2111, Q => 
                           registers_9_14_port);
   registers_reg_9_13_inst : DLH_X1 port map( G => n1992, D => n2114, Q => 
                           registers_9_13_port);
   registers_reg_9_12_inst : DLH_X1 port map( G => n1993, D => n2117, Q => 
                           registers_9_12_port);
   registers_reg_9_11_inst : DLH_X1 port map( G => n1992, D => n2120, Q => 
                           registers_9_11_port);
   registers_reg_9_10_inst : DLH_X1 port map( G => n1992, D => n2123, Q => 
                           registers_9_10_port);
   registers_reg_9_9_inst : DLH_X1 port map( G => n1992, D => n2126, Q => 
                           registers_9_9_port);
   registers_reg_9_8_inst : DLH_X1 port map( G => n1992, D => n2129, Q => 
                           registers_9_8_port);
   registers_reg_9_7_inst : DLH_X1 port map( G => n1992, D => n2132, Q => 
                           registers_9_7_port);
   registers_reg_9_6_inst : DLH_X1 port map( G => n1992, D => n2135, Q => 
                           registers_9_6_port);
   registers_reg_9_5_inst : DLH_X1 port map( G => n1992, D => n2138, Q => 
                           registers_9_5_port);
   registers_reg_9_4_inst : DLH_X1 port map( G => n1992, D => n2141, Q => 
                           registers_9_4_port);
   registers_reg_9_3_inst : DLH_X1 port map( G => n1992, D => n2144, Q => 
                           registers_9_3_port);
   registers_reg_9_2_inst : DLH_X1 port map( G => n1992, D => n2147, Q => 
                           registers_9_2_port);
   registers_reg_9_1_inst : DLH_X1 port map( G => n1993, D => n2150, Q => 
                           registers_9_1_port);
   registers_reg_9_0_inst : DLH_X1 port map( G => n1994, D => n2153, Q => 
                           registers_9_0_port);
   registers_reg_10_31_inst : DLH_X1 port map( G => n1997, D => n2059, Q => 
                           registers_10_31_port);
   registers_reg_10_30_inst : DLH_X1 port map( G => n1997, D => n2062, Q => 
                           registers_10_30_port);
   registers_reg_10_29_inst : DLH_X1 port map( G => n1997, D => n2065, Q => 
                           registers_10_29_port);
   registers_reg_10_28_inst : DLH_X1 port map( G => n1997, D => n2068, Q => 
                           registers_10_28_port);
   registers_reg_10_27_inst : DLH_X1 port map( G => n1997, D => n2071, Q => 
                           registers_10_27_port);
   registers_reg_10_26_inst : DLH_X1 port map( G => n1997, D => n2074, Q => 
                           registers_10_26_port);
   registers_reg_10_25_inst : DLH_X1 port map( G => n1997, D => n2077, Q => 
                           registers_10_25_port);
   registers_reg_10_24_inst : DLH_X1 port map( G => n1996, D => n2080, Q => 
                           registers_10_24_port);
   registers_reg_10_23_inst : DLH_X1 port map( G => n1996, D => n2083, Q => 
                           registers_10_23_port);
   registers_reg_10_22_inst : DLH_X1 port map( G => n1996, D => n2086, Q => 
                           registers_10_22_port);
   registers_reg_10_21_inst : DLH_X1 port map( G => n1996, D => n2089, Q => 
                           registers_10_21_port);
   registers_reg_10_20_inst : DLH_X1 port map( G => n1997, D => n2092, Q => 
                           registers_10_20_port);
   registers_reg_10_19_inst : DLH_X1 port map( G => n1996, D => n2095, Q => 
                           registers_10_19_port);
   registers_reg_10_18_inst : DLH_X1 port map( G => n1996, D => n2098, Q => 
                           registers_10_18_port);
   registers_reg_10_17_inst : DLH_X1 port map( G => n1997, D => n2101, Q => 
                           registers_10_17_port);
   registers_reg_10_16_inst : DLH_X1 port map( G => n1996, D => n2104, Q => 
                           registers_10_16_port);
   registers_reg_10_15_inst : DLH_X1 port map( G => n1996, D => n2107, Q => 
                           registers_10_15_port);
   registers_reg_10_14_inst : DLH_X1 port map( G => n1996, D => n2110, Q => 
                           registers_10_14_port);
   registers_reg_10_13_inst : DLH_X1 port map( G => n1995, D => n2113, Q => 
                           registers_10_13_port);
   registers_reg_10_12_inst : DLH_X1 port map( G => n1996, D => n2116, Q => 
                           registers_10_12_port);
   registers_reg_10_11_inst : DLH_X1 port map( G => n1995, D => n2119, Q => 
                           registers_10_11_port);
   registers_reg_10_10_inst : DLH_X1 port map( G => n1995, D => n2122, Q => 
                           registers_10_10_port);
   registers_reg_10_9_inst : DLH_X1 port map( G => n1995, D => n2125, Q => 
                           registers_10_9_port);
   registers_reg_10_8_inst : DLH_X1 port map( G => n1995, D => n2128, Q => 
                           registers_10_8_port);
   registers_reg_10_7_inst : DLH_X1 port map( G => n1995, D => n2131, Q => 
                           registers_10_7_port);
   registers_reg_10_6_inst : DLH_X1 port map( G => n1995, D => n2134, Q => 
                           registers_10_6_port);
   registers_reg_10_5_inst : DLH_X1 port map( G => n1995, D => n2137, Q => 
                           registers_10_5_port);
   registers_reg_10_4_inst : DLH_X1 port map( G => n1995, D => n2140, Q => 
                           registers_10_4_port);
   registers_reg_10_3_inst : DLH_X1 port map( G => n1995, D => n2143, Q => 
                           registers_10_3_port);
   registers_reg_10_2_inst : DLH_X1 port map( G => n1995, D => n2146, Q => 
                           registers_10_2_port);
   registers_reg_10_1_inst : DLH_X1 port map( G => n1996, D => n2149, Q => 
                           registers_10_1_port);
   registers_reg_10_0_inst : DLH_X1 port map( G => n1997, D => n2152, Q => 
                           registers_10_0_port);
   registers_reg_11_31_inst : DLH_X1 port map( G => n2000, D => n2059, Q => 
                           registers_11_31_port);
   registers_reg_11_30_inst : DLH_X1 port map( G => n2000, D => n2062, Q => 
                           registers_11_30_port);
   registers_reg_11_29_inst : DLH_X1 port map( G => n2000, D => n2065, Q => 
                           registers_11_29_port);
   registers_reg_11_28_inst : DLH_X1 port map( G => n2000, D => n2068, Q => 
                           registers_11_28_port);
   registers_reg_11_27_inst : DLH_X1 port map( G => n2000, D => n2071, Q => 
                           registers_11_27_port);
   registers_reg_11_26_inst : DLH_X1 port map( G => n2000, D => n2074, Q => 
                           registers_11_26_port);
   registers_reg_11_25_inst : DLH_X1 port map( G => n2000, D => n2077, Q => 
                           registers_11_25_port);
   registers_reg_11_24_inst : DLH_X1 port map( G => n1999, D => n2080, Q => 
                           registers_11_24_port);
   registers_reg_11_23_inst : DLH_X1 port map( G => n1999, D => n2083, Q => 
                           registers_11_23_port);
   registers_reg_11_22_inst : DLH_X1 port map( G => n1999, D => n2086, Q => 
                           registers_11_22_port);
   registers_reg_11_21_inst : DLH_X1 port map( G => n1999, D => n2089, Q => 
                           registers_11_21_port);
   registers_reg_11_20_inst : DLH_X1 port map( G => n2000, D => n2092, Q => 
                           registers_11_20_port);
   registers_reg_11_19_inst : DLH_X1 port map( G => n1999, D => n2095, Q => 
                           registers_11_19_port);
   registers_reg_11_18_inst : DLH_X1 port map( G => n1999, D => n2098, Q => 
                           registers_11_18_port);
   registers_reg_11_17_inst : DLH_X1 port map( G => n2000, D => n2101, Q => 
                           registers_11_17_port);
   registers_reg_11_16_inst : DLH_X1 port map( G => n1999, D => n2104, Q => 
                           registers_11_16_port);
   registers_reg_11_15_inst : DLH_X1 port map( G => n1999, D => n2107, Q => 
                           registers_11_15_port);
   registers_reg_11_14_inst : DLH_X1 port map( G => n1999, D => n2110, Q => 
                           registers_11_14_port);
   registers_reg_11_13_inst : DLH_X1 port map( G => n1998, D => n2113, Q => 
                           registers_11_13_port);
   registers_reg_11_12_inst : DLH_X1 port map( G => n1999, D => n2116, Q => 
                           registers_11_12_port);
   registers_reg_11_11_inst : DLH_X1 port map( G => n1998, D => n2119, Q => 
                           registers_11_11_port);
   registers_reg_11_10_inst : DLH_X1 port map( G => n1998, D => n2122, Q => 
                           registers_11_10_port);
   registers_reg_11_9_inst : DLH_X1 port map( G => n1998, D => n2125, Q => 
                           registers_11_9_port);
   registers_reg_11_8_inst : DLH_X1 port map( G => n1998, D => n2128, Q => 
                           registers_11_8_port);
   registers_reg_11_7_inst : DLH_X1 port map( G => n1998, D => n2131, Q => 
                           registers_11_7_port);
   registers_reg_11_6_inst : DLH_X1 port map( G => n1998, D => n2134, Q => 
                           registers_11_6_port);
   registers_reg_11_5_inst : DLH_X1 port map( G => n1998, D => n2137, Q => 
                           registers_11_5_port);
   registers_reg_11_4_inst : DLH_X1 port map( G => n1998, D => n2140, Q => 
                           registers_11_4_port);
   registers_reg_11_3_inst : DLH_X1 port map( G => n1998, D => n2143, Q => 
                           registers_11_3_port);
   registers_reg_11_2_inst : DLH_X1 port map( G => n1998, D => n2146, Q => 
                           registers_11_2_port);
   registers_reg_11_1_inst : DLH_X1 port map( G => n1999, D => n2149, Q => 
                           registers_11_1_port);
   registers_reg_11_0_inst : DLH_X1 port map( G => n2000, D => n2152, Q => 
                           registers_11_0_port);
   registers_reg_12_31_inst : DLH_X1 port map( G => n2001, D => n2059, Q => 
                           registers_12_31_port);
   registers_reg_12_30_inst : DLH_X1 port map( G => n2001, D => n2062, Q => 
                           registers_12_30_port);
   registers_reg_12_29_inst : DLH_X1 port map( G => n2001, D => n2065, Q => 
                           registers_12_29_port);
   registers_reg_12_28_inst : DLH_X1 port map( G => n2001, D => n2068, Q => 
                           registers_12_28_port);
   registers_reg_12_27_inst : DLH_X1 port map( G => n2001, D => n2071, Q => 
                           registers_12_27_port);
   registers_reg_12_26_inst : DLH_X1 port map( G => n2001, D => n2074, Q => 
                           registers_12_26_port);
   registers_reg_12_25_inst : DLH_X1 port map( G => n2001, D => n2077, Q => 
                           registers_12_25_port);
   registers_reg_12_24_inst : DLH_X1 port map( G => n2002, D => n2080, Q => 
                           registers_12_24_port);
   registers_reg_12_23_inst : DLH_X1 port map( G => n2002, D => n2083, Q => 
                           registers_12_23_port);
   registers_reg_12_22_inst : DLH_X1 port map( G => n2002, D => n2086, Q => 
                           registers_12_22_port);
   registers_reg_12_21_inst : DLH_X1 port map( G => n2002, D => n2089, Q => 
                           registers_12_21_port);
   registers_reg_12_20_inst : DLH_X1 port map( G => n2001, D => n2092, Q => 
                           registers_12_20_port);
   registers_reg_12_19_inst : DLH_X1 port map( G => n2002, D => n2095, Q => 
                           registers_12_19_port);
   registers_reg_12_18_inst : DLH_X1 port map( G => n2002, D => n2098, Q => 
                           registers_12_18_port);
   registers_reg_12_17_inst : DLH_X1 port map( G => n2001, D => n2101, Q => 
                           registers_12_17_port);
   registers_reg_12_16_inst : DLH_X1 port map( G => n2002, D => n2104, Q => 
                           registers_12_16_port);
   registers_reg_12_15_inst : DLH_X1 port map( G => n2002, D => n2107, Q => 
                           registers_12_15_port);
   registers_reg_12_14_inst : DLH_X1 port map( G => n2002, D => n2110, Q => 
                           registers_12_14_port);
   registers_reg_12_13_inst : DLH_X1 port map( G => n2002, D => n2113, Q => 
                           registers_12_13_port);
   registers_reg_12_12_inst : DLH_X1 port map( G => n2002, D => n2116, Q => 
                           registers_12_12_port);
   registers_reg_12_11_inst : DLH_X1 port map( G => n2003, D => n2119, Q => 
                           registers_12_11_port);
   registers_reg_12_10_inst : DLH_X1 port map( G => n2003, D => n2122, Q => 
                           registers_12_10_port);
   registers_reg_12_9_inst : DLH_X1 port map( G => n2003, D => n2125, Q => 
                           registers_12_9_port);
   registers_reg_12_8_inst : DLH_X1 port map( G => n2003, D => n2128, Q => 
                           registers_12_8_port);
   registers_reg_12_7_inst : DLH_X1 port map( G => n2003, D => n2131, Q => 
                           registers_12_7_port);
   registers_reg_12_6_inst : DLH_X1 port map( G => n2003, D => n2134, Q => 
                           registers_12_6_port);
   registers_reg_12_5_inst : DLH_X1 port map( G => n2003, D => n2137, Q => 
                           registers_12_5_port);
   registers_reg_12_4_inst : DLH_X1 port map( G => n2003, D => n2140, Q => 
                           registers_12_4_port);
   registers_reg_12_3_inst : DLH_X1 port map( G => n2003, D => n2143, Q => 
                           registers_12_3_port);
   registers_reg_12_2_inst : DLH_X1 port map( G => n2003, D => n2146, Q => 
                           registers_12_2_port);
   registers_reg_12_1_inst : DLH_X1 port map( G => n2001, D => n2149, Q => 
                           registers_12_1_port);
   registers_reg_12_0_inst : DLH_X1 port map( G => n2001, D => n2152, Q => 
                           registers_12_0_port);
   registers_reg_13_31_inst : DLH_X1 port map( G => n2004, D => n2059, Q => 
                           registers_13_31_port);
   registers_reg_13_30_inst : DLH_X1 port map( G => n2004, D => n2062, Q => 
                           registers_13_30_port);
   registers_reg_13_29_inst : DLH_X1 port map( G => n2004, D => n2065, Q => 
                           registers_13_29_port);
   registers_reg_13_28_inst : DLH_X1 port map( G => n2004, D => n2068, Q => 
                           registers_13_28_port);
   registers_reg_13_27_inst : DLH_X1 port map( G => n2004, D => n2071, Q => 
                           registers_13_27_port);
   registers_reg_13_26_inst : DLH_X1 port map( G => n2004, D => n2074, Q => 
                           registers_13_26_port);
   registers_reg_13_25_inst : DLH_X1 port map( G => n2004, D => n2077, Q => 
                           registers_13_25_port);
   registers_reg_13_24_inst : DLH_X1 port map( G => n2005, D => n2080, Q => 
                           registers_13_24_port);
   registers_reg_13_23_inst : DLH_X1 port map( G => n2005, D => n2083, Q => 
                           registers_13_23_port);
   registers_reg_13_22_inst : DLH_X1 port map( G => n2005, D => n2086, Q => 
                           registers_13_22_port);
   registers_reg_13_21_inst : DLH_X1 port map( G => n2005, D => n2089, Q => 
                           registers_13_21_port);
   registers_reg_13_20_inst : DLH_X1 port map( G => n2004, D => n2092, Q => 
                           registers_13_20_port);
   registers_reg_13_19_inst : DLH_X1 port map( G => n2005, D => n2095, Q => 
                           registers_13_19_port);
   registers_reg_13_18_inst : DLH_X1 port map( G => n2005, D => n2098, Q => 
                           registers_13_18_port);
   registers_reg_13_17_inst : DLH_X1 port map( G => n2004, D => n2101, Q => 
                           registers_13_17_port);
   registers_reg_13_16_inst : DLH_X1 port map( G => n2005, D => n2104, Q => 
                           registers_13_16_port);
   registers_reg_13_15_inst : DLH_X1 port map( G => n2005, D => n2107, Q => 
                           registers_13_15_port);
   registers_reg_13_14_inst : DLH_X1 port map( G => n2005, D => n2110, Q => 
                           registers_13_14_port);
   registers_reg_13_13_inst : DLH_X1 port map( G => n2005, D => n2113, Q => 
                           registers_13_13_port);
   registers_reg_13_12_inst : DLH_X1 port map( G => n2005, D => n2116, Q => 
                           registers_13_12_port);
   registers_reg_13_11_inst : DLH_X1 port map( G => n2006, D => n2119, Q => 
                           registers_13_11_port);
   registers_reg_13_10_inst : DLH_X1 port map( G => n2006, D => n2122, Q => 
                           registers_13_10_port);
   registers_reg_13_9_inst : DLH_X1 port map( G => n2006, D => n2125, Q => 
                           registers_13_9_port);
   registers_reg_13_8_inst : DLH_X1 port map( G => n2006, D => n2128, Q => 
                           registers_13_8_port);
   registers_reg_13_7_inst : DLH_X1 port map( G => n2006, D => n2131, Q => 
                           registers_13_7_port);
   registers_reg_13_6_inst : DLH_X1 port map( G => n2006, D => n2134, Q => 
                           registers_13_6_port);
   registers_reg_13_5_inst : DLH_X1 port map( G => n2006, D => n2137, Q => 
                           registers_13_5_port);
   registers_reg_13_4_inst : DLH_X1 port map( G => n2006, D => n2140, Q => 
                           registers_13_4_port);
   registers_reg_13_3_inst : DLH_X1 port map( G => n2006, D => n2143, Q => 
                           registers_13_3_port);
   registers_reg_13_2_inst : DLH_X1 port map( G => n2006, D => n2146, Q => 
                           registers_13_2_port);
   registers_reg_13_1_inst : DLH_X1 port map( G => n2004, D => n2149, Q => 
                           registers_13_1_port);
   registers_reg_13_0_inst : DLH_X1 port map( G => n2004, D => n2152, Q => 
                           registers_13_0_port);
   registers_reg_14_31_inst : DLH_X1 port map( G => n2007, D => n2059, Q => 
                           registers_14_31_port);
   registers_reg_14_30_inst : DLH_X1 port map( G => n2007, D => n2062, Q => 
                           registers_14_30_port);
   registers_reg_14_29_inst : DLH_X1 port map( G => n2007, D => n2065, Q => 
                           registers_14_29_port);
   registers_reg_14_28_inst : DLH_X1 port map( G => n2007, D => n2068, Q => 
                           registers_14_28_port);
   registers_reg_14_27_inst : DLH_X1 port map( G => n2007, D => n2071, Q => 
                           registers_14_27_port);
   registers_reg_14_26_inst : DLH_X1 port map( G => n2007, D => n2074, Q => 
                           registers_14_26_port);
   registers_reg_14_25_inst : DLH_X1 port map( G => n2007, D => n2077, Q => 
                           registers_14_25_port);
   registers_reg_14_24_inst : DLH_X1 port map( G => n2008, D => n2080, Q => 
                           registers_14_24_port);
   registers_reg_14_23_inst : DLH_X1 port map( G => n2008, D => n2083, Q => 
                           registers_14_23_port);
   registers_reg_14_22_inst : DLH_X1 port map( G => n2008, D => n2086, Q => 
                           registers_14_22_port);
   registers_reg_14_21_inst : DLH_X1 port map( G => n2008, D => n2089, Q => 
                           registers_14_21_port);
   registers_reg_14_20_inst : DLH_X1 port map( G => n2007, D => n2092, Q => 
                           registers_14_20_port);
   registers_reg_14_19_inst : DLH_X1 port map( G => n2008, D => n2095, Q => 
                           registers_14_19_port);
   registers_reg_14_18_inst : DLH_X1 port map( G => n2008, D => n2098, Q => 
                           registers_14_18_port);
   registers_reg_14_17_inst : DLH_X1 port map( G => n2007, D => n2101, Q => 
                           registers_14_17_port);
   registers_reg_14_16_inst : DLH_X1 port map( G => n2008, D => n2104, Q => 
                           registers_14_16_port);
   registers_reg_14_15_inst : DLH_X1 port map( G => n2008, D => n2107, Q => 
                           registers_14_15_port);
   registers_reg_14_14_inst : DLH_X1 port map( G => n2008, D => n2110, Q => 
                           registers_14_14_port);
   registers_reg_14_13_inst : DLH_X1 port map( G => n2008, D => n2113, Q => 
                           registers_14_13_port);
   registers_reg_14_12_inst : DLH_X1 port map( G => n2008, D => n2116, Q => 
                           registers_14_12_port);
   registers_reg_14_11_inst : DLH_X1 port map( G => n2009, D => n2119, Q => 
                           registers_14_11_port);
   registers_reg_14_10_inst : DLH_X1 port map( G => n2009, D => n2122, Q => 
                           registers_14_10_port);
   registers_reg_14_9_inst : DLH_X1 port map( G => n2009, D => n2125, Q => 
                           registers_14_9_port);
   registers_reg_14_8_inst : DLH_X1 port map( G => n2009, D => n2128, Q => 
                           registers_14_8_port);
   registers_reg_14_7_inst : DLH_X1 port map( G => n2009, D => n2131, Q => 
                           registers_14_7_port);
   registers_reg_14_6_inst : DLH_X1 port map( G => n2009, D => n2134, Q => 
                           registers_14_6_port);
   registers_reg_14_5_inst : DLH_X1 port map( G => n2009, D => n2137, Q => 
                           registers_14_5_port);
   registers_reg_14_4_inst : DLH_X1 port map( G => n2009, D => n2140, Q => 
                           registers_14_4_port);
   registers_reg_14_3_inst : DLH_X1 port map( G => n2009, D => n2143, Q => 
                           registers_14_3_port);
   registers_reg_14_2_inst : DLH_X1 port map( G => n2009, D => n2146, Q => 
                           registers_14_2_port);
   registers_reg_14_1_inst : DLH_X1 port map( G => n2007, D => n2149, Q => 
                           registers_14_1_port);
   registers_reg_14_0_inst : DLH_X1 port map( G => n2007, D => n2152, Q => 
                           registers_14_0_port);
   registers_reg_15_31_inst : DLH_X1 port map( G => n2010, D => n2059, Q => 
                           registers_15_31_port);
   registers_reg_15_30_inst : DLH_X1 port map( G => n2010, D => n2062, Q => 
                           registers_15_30_port);
   registers_reg_15_29_inst : DLH_X1 port map( G => n2010, D => n2065, Q => 
                           registers_15_29_port);
   registers_reg_15_28_inst : DLH_X1 port map( G => n2010, D => n2068, Q => 
                           registers_15_28_port);
   registers_reg_15_27_inst : DLH_X1 port map( G => n2010, D => n2071, Q => 
                           registers_15_27_port);
   registers_reg_15_26_inst : DLH_X1 port map( G => n2010, D => n2074, Q => 
                           registers_15_26_port);
   registers_reg_15_25_inst : DLH_X1 port map( G => n2010, D => n2077, Q => 
                           registers_15_25_port);
   registers_reg_15_24_inst : DLH_X1 port map( G => n2011, D => n2080, Q => 
                           registers_15_24_port);
   registers_reg_15_23_inst : DLH_X1 port map( G => n2011, D => n2083, Q => 
                           registers_15_23_port);
   registers_reg_15_22_inst : DLH_X1 port map( G => n2011, D => n2086, Q => 
                           registers_15_22_port);
   registers_reg_15_21_inst : DLH_X1 port map( G => n2011, D => n2089, Q => 
                           registers_15_21_port);
   registers_reg_15_20_inst : DLH_X1 port map( G => n2010, D => n2092, Q => 
                           registers_15_20_port);
   registers_reg_15_19_inst : DLH_X1 port map( G => n2011, D => n2095, Q => 
                           registers_15_19_port);
   registers_reg_15_18_inst : DLH_X1 port map( G => n2011, D => n2098, Q => 
                           registers_15_18_port);
   registers_reg_15_17_inst : DLH_X1 port map( G => n2010, D => n2101, Q => 
                           registers_15_17_port);
   registers_reg_15_16_inst : DLH_X1 port map( G => n2011, D => n2104, Q => 
                           registers_15_16_port);
   registers_reg_15_15_inst : DLH_X1 port map( G => n2011, D => n2107, Q => 
                           registers_15_15_port);
   registers_reg_15_14_inst : DLH_X1 port map( G => n2011, D => n2110, Q => 
                           registers_15_14_port);
   registers_reg_15_13_inst : DLH_X1 port map( G => n2011, D => n2113, Q => 
                           registers_15_13_port);
   registers_reg_15_12_inst : DLH_X1 port map( G => n2011, D => n2116, Q => 
                           registers_15_12_port);
   registers_reg_15_11_inst : DLH_X1 port map( G => n2012, D => n2119, Q => 
                           registers_15_11_port);
   registers_reg_15_10_inst : DLH_X1 port map( G => n2012, D => n2122, Q => 
                           registers_15_10_port);
   registers_reg_15_9_inst : DLH_X1 port map( G => n2012, D => n2125, Q => 
                           registers_15_9_port);
   registers_reg_15_8_inst : DLH_X1 port map( G => n2012, D => n2128, Q => 
                           registers_15_8_port);
   registers_reg_15_7_inst : DLH_X1 port map( G => n2012, D => n2131, Q => 
                           registers_15_7_port);
   registers_reg_15_6_inst : DLH_X1 port map( G => n2012, D => n2134, Q => 
                           registers_15_6_port);
   registers_reg_15_5_inst : DLH_X1 port map( G => n2012, D => n2137, Q => 
                           registers_15_5_port);
   registers_reg_15_4_inst : DLH_X1 port map( G => n2012, D => n2140, Q => 
                           registers_15_4_port);
   registers_reg_15_3_inst : DLH_X1 port map( G => n2012, D => n2143, Q => 
                           registers_15_3_port);
   registers_reg_15_2_inst : DLH_X1 port map( G => n2012, D => n2146, Q => 
                           registers_15_2_port);
   registers_reg_15_1_inst : DLH_X1 port map( G => n2010, D => n2149, Q => 
                           registers_15_1_port);
   registers_reg_15_0_inst : DLH_X1 port map( G => n2010, D => n2152, Q => 
                           registers_15_0_port);
   registers_reg_16_31_inst : DLH_X1 port map( G => n2013, D => n2059, Q => 
                           registers_16_31_port);
   registers_reg_16_30_inst : DLH_X1 port map( G => n2013, D => n2062, Q => 
                           registers_16_30_port);
   registers_reg_16_29_inst : DLH_X1 port map( G => n2013, D => n2065, Q => 
                           registers_16_29_port);
   registers_reg_16_28_inst : DLH_X1 port map( G => n2013, D => n2068, Q => 
                           registers_16_28_port);
   registers_reg_16_27_inst : DLH_X1 port map( G => n2013, D => n2071, Q => 
                           registers_16_27_port);
   registers_reg_16_26_inst : DLH_X1 port map( G => n2013, D => n2074, Q => 
                           registers_16_26_port);
   registers_reg_16_25_inst : DLH_X1 port map( G => n2013, D => n2077, Q => 
                           registers_16_25_port);
   registers_reg_16_24_inst : DLH_X1 port map( G => n2014, D => n2080, Q => 
                           registers_16_24_port);
   registers_reg_16_23_inst : DLH_X1 port map( G => n2014, D => n2083, Q => 
                           registers_16_23_port);
   registers_reg_16_22_inst : DLH_X1 port map( G => n2014, D => n2086, Q => 
                           registers_16_22_port);
   registers_reg_16_21_inst : DLH_X1 port map( G => n2014, D => n2089, Q => 
                           registers_16_21_port);
   registers_reg_16_20_inst : DLH_X1 port map( G => n2013, D => n2092, Q => 
                           registers_16_20_port);
   registers_reg_16_19_inst : DLH_X1 port map( G => n2014, D => n2095, Q => 
                           registers_16_19_port);
   registers_reg_16_18_inst : DLH_X1 port map( G => n2014, D => n2098, Q => 
                           registers_16_18_port);
   registers_reg_16_17_inst : DLH_X1 port map( G => n2013, D => n2101, Q => 
                           registers_16_17_port);
   registers_reg_16_16_inst : DLH_X1 port map( G => n2014, D => n2104, Q => 
                           registers_16_16_port);
   registers_reg_16_15_inst : DLH_X1 port map( G => n2014, D => n2107, Q => 
                           registers_16_15_port);
   registers_reg_16_14_inst : DLH_X1 port map( G => n2014, D => n2110, Q => 
                           registers_16_14_port);
   registers_reg_16_13_inst : DLH_X1 port map( G => n2014, D => n2113, Q => 
                           registers_16_13_port);
   registers_reg_16_12_inst : DLH_X1 port map( G => n2014, D => n2116, Q => 
                           registers_16_12_port);
   registers_reg_16_11_inst : DLH_X1 port map( G => n2015, D => n2119, Q => 
                           registers_16_11_port);
   registers_reg_16_10_inst : DLH_X1 port map( G => n2015, D => n2122, Q => 
                           registers_16_10_port);
   registers_reg_16_9_inst : DLH_X1 port map( G => n2015, D => n2125, Q => 
                           registers_16_9_port);
   registers_reg_16_8_inst : DLH_X1 port map( G => n2015, D => n2128, Q => 
                           registers_16_8_port);
   registers_reg_16_7_inst : DLH_X1 port map( G => n2015, D => n2131, Q => 
                           registers_16_7_port);
   registers_reg_16_6_inst : DLH_X1 port map( G => n2015, D => n2134, Q => 
                           registers_16_6_port);
   registers_reg_16_5_inst : DLH_X1 port map( G => n2015, D => n2137, Q => 
                           registers_16_5_port);
   registers_reg_16_4_inst : DLH_X1 port map( G => n2015, D => n2140, Q => 
                           registers_16_4_port);
   registers_reg_16_3_inst : DLH_X1 port map( G => n2015, D => n2143, Q => 
                           registers_16_3_port);
   registers_reg_16_2_inst : DLH_X1 port map( G => n2015, D => n2146, Q => 
                           registers_16_2_port);
   registers_reg_16_1_inst : DLH_X1 port map( G => n2013, D => n2149, Q => 
                           registers_16_1_port);
   registers_reg_16_0_inst : DLH_X1 port map( G => n2013, D => n2152, Q => 
                           registers_16_0_port);
   registers_reg_17_31_inst : DLH_X1 port map( G => n2016, D => n2059, Q => 
                           registers_17_31_port);
   registers_reg_17_30_inst : DLH_X1 port map( G => n2016, D => n2062, Q => 
                           registers_17_30_port);
   registers_reg_17_29_inst : DLH_X1 port map( G => n2016, D => n2065, Q => 
                           registers_17_29_port);
   registers_reg_17_28_inst : DLH_X1 port map( G => n2016, D => n2068, Q => 
                           registers_17_28_port);
   registers_reg_17_27_inst : DLH_X1 port map( G => n2016, D => n2071, Q => 
                           registers_17_27_port);
   registers_reg_17_26_inst : DLH_X1 port map( G => n2016, D => n2074, Q => 
                           registers_17_26_port);
   registers_reg_17_25_inst : DLH_X1 port map( G => n2016, D => n2077, Q => 
                           registers_17_25_port);
   registers_reg_17_24_inst : DLH_X1 port map( G => n2017, D => n2080, Q => 
                           registers_17_24_port);
   registers_reg_17_23_inst : DLH_X1 port map( G => n2017, D => n2083, Q => 
                           registers_17_23_port);
   registers_reg_17_22_inst : DLH_X1 port map( G => n2017, D => n2086, Q => 
                           registers_17_22_port);
   registers_reg_17_21_inst : DLH_X1 port map( G => n2017, D => n2089, Q => 
                           registers_17_21_port);
   registers_reg_17_20_inst : DLH_X1 port map( G => n2016, D => n2092, Q => 
                           registers_17_20_port);
   registers_reg_17_19_inst : DLH_X1 port map( G => n2017, D => n2095, Q => 
                           registers_17_19_port);
   registers_reg_17_18_inst : DLH_X1 port map( G => n2017, D => n2098, Q => 
                           registers_17_18_port);
   registers_reg_17_17_inst : DLH_X1 port map( G => n2016, D => n2101, Q => 
                           registers_17_17_port);
   registers_reg_17_16_inst : DLH_X1 port map( G => n2017, D => n2104, Q => 
                           registers_17_16_port);
   registers_reg_17_15_inst : DLH_X1 port map( G => n2017, D => n2107, Q => 
                           registers_17_15_port);
   registers_reg_17_14_inst : DLH_X1 port map( G => n2017, D => n2110, Q => 
                           registers_17_14_port);
   registers_reg_17_13_inst : DLH_X1 port map( G => n2017, D => n2113, Q => 
                           registers_17_13_port);
   registers_reg_17_12_inst : DLH_X1 port map( G => n2017, D => n2116, Q => 
                           registers_17_12_port);
   registers_reg_17_11_inst : DLH_X1 port map( G => n2018, D => n2119, Q => 
                           registers_17_11_port);
   registers_reg_17_10_inst : DLH_X1 port map( G => n2018, D => n2122, Q => 
                           registers_17_10_port);
   registers_reg_17_9_inst : DLH_X1 port map( G => n2018, D => n2125, Q => 
                           registers_17_9_port);
   registers_reg_17_8_inst : DLH_X1 port map( G => n2018, D => n2128, Q => 
                           registers_17_8_port);
   registers_reg_17_7_inst : DLH_X1 port map( G => n2018, D => n2131, Q => 
                           registers_17_7_port);
   registers_reg_17_6_inst : DLH_X1 port map( G => n2018, D => n2134, Q => 
                           registers_17_6_port);
   registers_reg_17_5_inst : DLH_X1 port map( G => n2018, D => n2137, Q => 
                           registers_17_5_port);
   registers_reg_17_4_inst : DLH_X1 port map( G => n2018, D => n2140, Q => 
                           registers_17_4_port);
   registers_reg_17_3_inst : DLH_X1 port map( G => n2018, D => n2143, Q => 
                           registers_17_3_port);
   registers_reg_17_2_inst : DLH_X1 port map( G => n2018, D => n2146, Q => 
                           registers_17_2_port);
   registers_reg_17_1_inst : DLH_X1 port map( G => n2016, D => n2149, Q => 
                           registers_17_1_port);
   registers_reg_17_0_inst : DLH_X1 port map( G => n2016, D => n2152, Q => 
                           registers_17_0_port);
   registers_reg_18_31_inst : DLH_X1 port map( G => n2019, D => n2059, Q => 
                           registers_18_31_port);
   registers_reg_18_30_inst : DLH_X1 port map( G => n2019, D => n2062, Q => 
                           registers_18_30_port);
   registers_reg_18_29_inst : DLH_X1 port map( G => n2019, D => n2065, Q => 
                           registers_18_29_port);
   registers_reg_18_28_inst : DLH_X1 port map( G => n2019, D => n2068, Q => 
                           registers_18_28_port);
   registers_reg_18_27_inst : DLH_X1 port map( G => n2019, D => n2071, Q => 
                           registers_18_27_port);
   registers_reg_18_26_inst : DLH_X1 port map( G => n2019, D => n2074, Q => 
                           registers_18_26_port);
   registers_reg_18_25_inst : DLH_X1 port map( G => n2019, D => n2077, Q => 
                           registers_18_25_port);
   registers_reg_18_24_inst : DLH_X1 port map( G => n2020, D => n2080, Q => 
                           registers_18_24_port);
   registers_reg_18_23_inst : DLH_X1 port map( G => n2020, D => n2083, Q => 
                           registers_18_23_port);
   registers_reg_18_22_inst : DLH_X1 port map( G => n2020, D => n2086, Q => 
                           registers_18_22_port);
   registers_reg_18_21_inst : DLH_X1 port map( G => n2020, D => n2089, Q => 
                           registers_18_21_port);
   registers_reg_18_20_inst : DLH_X1 port map( G => n2019, D => n2092, Q => 
                           registers_18_20_port);
   registers_reg_18_19_inst : DLH_X1 port map( G => n2020, D => n2095, Q => 
                           registers_18_19_port);
   registers_reg_18_18_inst : DLH_X1 port map( G => n2020, D => n2098, Q => 
                           registers_18_18_port);
   registers_reg_18_17_inst : DLH_X1 port map( G => n2019, D => n2101, Q => 
                           registers_18_17_port);
   registers_reg_18_16_inst : DLH_X1 port map( G => n2020, D => n2104, Q => 
                           registers_18_16_port);
   registers_reg_18_15_inst : DLH_X1 port map( G => n2020, D => n2107, Q => 
                           registers_18_15_port);
   registers_reg_18_14_inst : DLH_X1 port map( G => n2020, D => n2110, Q => 
                           registers_18_14_port);
   registers_reg_18_13_inst : DLH_X1 port map( G => n2020, D => n2113, Q => 
                           registers_18_13_port);
   registers_reg_18_12_inst : DLH_X1 port map( G => n2020, D => n2116, Q => 
                           registers_18_12_port);
   registers_reg_18_11_inst : DLH_X1 port map( G => n2021, D => n2119, Q => 
                           registers_18_11_port);
   registers_reg_18_10_inst : DLH_X1 port map( G => n2021, D => n2122, Q => 
                           registers_18_10_port);
   registers_reg_18_9_inst : DLH_X1 port map( G => n2021, D => n2125, Q => 
                           registers_18_9_port);
   registers_reg_18_8_inst : DLH_X1 port map( G => n2021, D => n2128, Q => 
                           registers_18_8_port);
   registers_reg_18_7_inst : DLH_X1 port map( G => n2021, D => n2131, Q => 
                           registers_18_7_port);
   registers_reg_18_6_inst : DLH_X1 port map( G => n2021, D => n2134, Q => 
                           registers_18_6_port);
   registers_reg_18_5_inst : DLH_X1 port map( G => n2021, D => n2137, Q => 
                           registers_18_5_port);
   registers_reg_18_4_inst : DLH_X1 port map( G => n2021, D => n2140, Q => 
                           registers_18_4_port);
   registers_reg_18_3_inst : DLH_X1 port map( G => n2021, D => n2143, Q => 
                           registers_18_3_port);
   registers_reg_18_2_inst : DLH_X1 port map( G => n2021, D => n2146, Q => 
                           registers_18_2_port);
   registers_reg_18_1_inst : DLH_X1 port map( G => n2019, D => n2149, Q => 
                           registers_18_1_port);
   registers_reg_18_0_inst : DLH_X1 port map( G => n2019, D => n2152, Q => 
                           registers_18_0_port);
   registers_reg_19_31_inst : DLH_X1 port map( G => n2022, D => n2059, Q => 
                           registers_19_31_port);
   registers_reg_19_30_inst : DLH_X1 port map( G => n2022, D => n2062, Q => 
                           registers_19_30_port);
   registers_reg_19_29_inst : DLH_X1 port map( G => n2022, D => n2065, Q => 
                           registers_19_29_port);
   registers_reg_19_28_inst : DLH_X1 port map( G => n2022, D => n2068, Q => 
                           registers_19_28_port);
   registers_reg_19_27_inst : DLH_X1 port map( G => n2022, D => n2071, Q => 
                           registers_19_27_port);
   registers_reg_19_26_inst : DLH_X1 port map( G => n2022, D => n2074, Q => 
                           registers_19_26_port);
   registers_reg_19_25_inst : DLH_X1 port map( G => n2022, D => n2077, Q => 
                           registers_19_25_port);
   registers_reg_19_24_inst : DLH_X1 port map( G => n2023, D => n2080, Q => 
                           registers_19_24_port);
   registers_reg_19_23_inst : DLH_X1 port map( G => n2023, D => n2083, Q => 
                           registers_19_23_port);
   registers_reg_19_22_inst : DLH_X1 port map( G => n2023, D => n2086, Q => 
                           registers_19_22_port);
   registers_reg_19_21_inst : DLH_X1 port map( G => n2023, D => n2089, Q => 
                           registers_19_21_port);
   registers_reg_19_20_inst : DLH_X1 port map( G => n2022, D => n2092, Q => 
                           registers_19_20_port);
   registers_reg_19_19_inst : DLH_X1 port map( G => n2023, D => n2095, Q => 
                           registers_19_19_port);
   registers_reg_19_18_inst : DLH_X1 port map( G => n2023, D => n2098, Q => 
                           registers_19_18_port);
   registers_reg_19_17_inst : DLH_X1 port map( G => n2022, D => n2101, Q => 
                           registers_19_17_port);
   registers_reg_19_16_inst : DLH_X1 port map( G => n2023, D => n2104, Q => 
                           registers_19_16_port);
   registers_reg_19_15_inst : DLH_X1 port map( G => n2023, D => n2107, Q => 
                           registers_19_15_port);
   registers_reg_19_14_inst : DLH_X1 port map( G => n2023, D => n2110, Q => 
                           registers_19_14_port);
   registers_reg_19_13_inst : DLH_X1 port map( G => n2023, D => n2113, Q => 
                           registers_19_13_port);
   registers_reg_19_12_inst : DLH_X1 port map( G => n2023, D => n2116, Q => 
                           registers_19_12_port);
   registers_reg_19_11_inst : DLH_X1 port map( G => n2024, D => n2119, Q => 
                           registers_19_11_port);
   registers_reg_19_10_inst : DLH_X1 port map( G => n2024, D => n2122, Q => 
                           registers_19_10_port);
   registers_reg_19_9_inst : DLH_X1 port map( G => n2024, D => n2125, Q => 
                           registers_19_9_port);
   registers_reg_19_8_inst : DLH_X1 port map( G => n2024, D => n2128, Q => 
                           registers_19_8_port);
   registers_reg_19_7_inst : DLH_X1 port map( G => n2024, D => n2131, Q => 
                           registers_19_7_port);
   registers_reg_19_6_inst : DLH_X1 port map( G => n2024, D => n2134, Q => 
                           registers_19_6_port);
   registers_reg_19_5_inst : DLH_X1 port map( G => n2024, D => n2137, Q => 
                           registers_19_5_port);
   registers_reg_19_4_inst : DLH_X1 port map( G => n2024, D => n2140, Q => 
                           registers_19_4_port);
   registers_reg_19_3_inst : DLH_X1 port map( G => n2024, D => n2143, Q => 
                           registers_19_3_port);
   registers_reg_19_2_inst : DLH_X1 port map( G => n2024, D => n2146, Q => 
                           registers_19_2_port);
   registers_reg_19_1_inst : DLH_X1 port map( G => n2022, D => n2149, Q => 
                           registers_19_1_port);
   registers_reg_19_0_inst : DLH_X1 port map( G => n2022, D => n2152, Q => 
                           registers_19_0_port);
   registers_reg_20_31_inst : DLH_X1 port map( G => n2025, D => n2059, Q => 
                           registers_20_31_port);
   registers_reg_20_30_inst : DLH_X1 port map( G => n2025, D => n2062, Q => 
                           registers_20_30_port);
   registers_reg_20_29_inst : DLH_X1 port map( G => n2025, D => n2065, Q => 
                           registers_20_29_port);
   registers_reg_20_28_inst : DLH_X1 port map( G => n2025, D => n2068, Q => 
                           registers_20_28_port);
   registers_reg_20_27_inst : DLH_X1 port map( G => n2025, D => n2071, Q => 
                           registers_20_27_port);
   registers_reg_20_26_inst : DLH_X1 port map( G => n2025, D => n2074, Q => 
                           registers_20_26_port);
   registers_reg_20_25_inst : DLH_X1 port map( G => n2025, D => n2077, Q => 
                           registers_20_25_port);
   registers_reg_20_24_inst : DLH_X1 port map( G => n2026, D => n2080, Q => 
                           registers_20_24_port);
   registers_reg_20_23_inst : DLH_X1 port map( G => n2026, D => n2083, Q => 
                           registers_20_23_port);
   registers_reg_20_22_inst : DLH_X1 port map( G => n2026, D => n2086, Q => 
                           registers_20_22_port);
   registers_reg_20_21_inst : DLH_X1 port map( G => n2026, D => n2089, Q => 
                           registers_20_21_port);
   registers_reg_20_20_inst : DLH_X1 port map( G => n2025, D => n2092, Q => 
                           registers_20_20_port);
   registers_reg_20_19_inst : DLH_X1 port map( G => n2026, D => n2095, Q => 
                           registers_20_19_port);
   registers_reg_20_18_inst : DLH_X1 port map( G => n2026, D => n2098, Q => 
                           registers_20_18_port);
   registers_reg_20_17_inst : DLH_X1 port map( G => n2025, D => n2101, Q => 
                           registers_20_17_port);
   registers_reg_20_16_inst : DLH_X1 port map( G => n2026, D => n2104, Q => 
                           registers_20_16_port);
   registers_reg_20_15_inst : DLH_X1 port map( G => n2026, D => n2107, Q => 
                           registers_20_15_port);
   registers_reg_20_14_inst : DLH_X1 port map( G => n2026, D => n2110, Q => 
                           registers_20_14_port);
   registers_reg_20_13_inst : DLH_X1 port map( G => n2026, D => n2113, Q => 
                           registers_20_13_port);
   registers_reg_20_12_inst : DLH_X1 port map( G => n2026, D => n2116, Q => 
                           registers_20_12_port);
   registers_reg_20_11_inst : DLH_X1 port map( G => n2027, D => n2119, Q => 
                           registers_20_11_port);
   registers_reg_20_10_inst : DLH_X1 port map( G => n2027, D => n2122, Q => 
                           registers_20_10_port);
   registers_reg_20_9_inst : DLH_X1 port map( G => n2027, D => n2125, Q => 
                           registers_20_9_port);
   registers_reg_20_8_inst : DLH_X1 port map( G => n2027, D => n2128, Q => 
                           registers_20_8_port);
   registers_reg_20_7_inst : DLH_X1 port map( G => n2027, D => n2131, Q => 
                           registers_20_7_port);
   registers_reg_20_6_inst : DLH_X1 port map( G => n2027, D => n2134, Q => 
                           registers_20_6_port);
   registers_reg_20_5_inst : DLH_X1 port map( G => n2027, D => n2137, Q => 
                           registers_20_5_port);
   registers_reg_20_4_inst : DLH_X1 port map( G => n2027, D => n2140, Q => 
                           registers_20_4_port);
   registers_reg_20_3_inst : DLH_X1 port map( G => n2027, D => n2143, Q => 
                           registers_20_3_port);
   registers_reg_20_2_inst : DLH_X1 port map( G => n2027, D => n2146, Q => 
                           registers_20_2_port);
   registers_reg_20_1_inst : DLH_X1 port map( G => n2025, D => n2149, Q => 
                           registers_20_1_port);
   registers_reg_20_0_inst : DLH_X1 port map( G => n2025, D => n2152, Q => 
                           registers_20_0_port);
   registers_reg_21_31_inst : DLH_X1 port map( G => n2028, D => n2058, Q => 
                           registers_21_31_port);
   registers_reg_21_30_inst : DLH_X1 port map( G => n2028, D => n2061, Q => 
                           registers_21_30_port);
   registers_reg_21_29_inst : DLH_X1 port map( G => n2028, D => n2064, Q => 
                           registers_21_29_port);
   registers_reg_21_28_inst : DLH_X1 port map( G => n2028, D => n2067, Q => 
                           registers_21_28_port);
   registers_reg_21_27_inst : DLH_X1 port map( G => n2028, D => n2070, Q => 
                           registers_21_27_port);
   registers_reg_21_26_inst : DLH_X1 port map( G => n2028, D => n2073, Q => 
                           registers_21_26_port);
   registers_reg_21_25_inst : DLH_X1 port map( G => n2028, D => n2076, Q => 
                           registers_21_25_port);
   registers_reg_21_24_inst : DLH_X1 port map( G => n2029, D => n2079, Q => 
                           registers_21_24_port);
   registers_reg_21_23_inst : DLH_X1 port map( G => n2029, D => n2082, Q => 
                           registers_21_23_port);
   registers_reg_21_22_inst : DLH_X1 port map( G => n2029, D => n2085, Q => 
                           registers_21_22_port);
   registers_reg_21_21_inst : DLH_X1 port map( G => n2029, D => n2088, Q => 
                           registers_21_21_port);
   registers_reg_21_20_inst : DLH_X1 port map( G => n2028, D => n2091, Q => 
                           registers_21_20_port);
   registers_reg_21_19_inst : DLH_X1 port map( G => n2029, D => n2094, Q => 
                           registers_21_19_port);
   registers_reg_21_18_inst : DLH_X1 port map( G => n2029, D => n2097, Q => 
                           registers_21_18_port);
   registers_reg_21_17_inst : DLH_X1 port map( G => n2028, D => n2100, Q => 
                           registers_21_17_port);
   registers_reg_21_16_inst : DLH_X1 port map( G => n2029, D => n2103, Q => 
                           registers_21_16_port);
   registers_reg_21_15_inst : DLH_X1 port map( G => n2029, D => n2106, Q => 
                           registers_21_15_port);
   registers_reg_21_14_inst : DLH_X1 port map( G => n2029, D => n2109, Q => 
                           registers_21_14_port);
   registers_reg_21_13_inst : DLH_X1 port map( G => n2029, D => n2112, Q => 
                           registers_21_13_port);
   registers_reg_21_12_inst : DLH_X1 port map( G => n2029, D => n2115, Q => 
                           registers_21_12_port);
   registers_reg_21_11_inst : DLH_X1 port map( G => n2030, D => n2118, Q => 
                           registers_21_11_port);
   registers_reg_21_10_inst : DLH_X1 port map( G => n2030, D => n2121, Q => 
                           registers_21_10_port);
   registers_reg_21_9_inst : DLH_X1 port map( G => n2030, D => n2124, Q => 
                           registers_21_9_port);
   registers_reg_21_8_inst : DLH_X1 port map( G => n2030, D => n2127, Q => 
                           registers_21_8_port);
   registers_reg_21_7_inst : DLH_X1 port map( G => n2030, D => n2130, Q => 
                           registers_21_7_port);
   registers_reg_21_6_inst : DLH_X1 port map( G => n2030, D => n2133, Q => 
                           registers_21_6_port);
   registers_reg_21_5_inst : DLH_X1 port map( G => n2030, D => n2136, Q => 
                           registers_21_5_port);
   registers_reg_21_4_inst : DLH_X1 port map( G => n2030, D => n2139, Q => 
                           registers_21_4_port);
   registers_reg_21_3_inst : DLH_X1 port map( G => n2030, D => n2142, Q => 
                           registers_21_3_port);
   registers_reg_21_2_inst : DLH_X1 port map( G => n2030, D => n2145, Q => 
                           registers_21_2_port);
   registers_reg_21_1_inst : DLH_X1 port map( G => n2028, D => n2148, Q => 
                           registers_21_1_port);
   registers_reg_21_0_inst : DLH_X1 port map( G => n2028, D => n2151, Q => 
                           registers_21_0_port);
   registers_reg_22_31_inst : DLH_X1 port map( G => n2031, D => n2058, Q => 
                           registers_22_31_port);
   registers_reg_22_30_inst : DLH_X1 port map( G => n2031, D => n2061, Q => 
                           registers_22_30_port);
   registers_reg_22_29_inst : DLH_X1 port map( G => n2031, D => n2064, Q => 
                           registers_22_29_port);
   registers_reg_22_28_inst : DLH_X1 port map( G => n2031, D => n2067, Q => 
                           registers_22_28_port);
   registers_reg_22_27_inst : DLH_X1 port map( G => n2031, D => n2070, Q => 
                           registers_22_27_port);
   registers_reg_22_26_inst : DLH_X1 port map( G => n2031, D => n2073, Q => 
                           registers_22_26_port);
   registers_reg_22_25_inst : DLH_X1 port map( G => n2031, D => n2076, Q => 
                           registers_22_25_port);
   registers_reg_22_24_inst : DLH_X1 port map( G => n2032, D => n2079, Q => 
                           registers_22_24_port);
   registers_reg_22_23_inst : DLH_X1 port map( G => n2032, D => n2082, Q => 
                           registers_22_23_port);
   registers_reg_22_22_inst : DLH_X1 port map( G => n2032, D => n2085, Q => 
                           registers_22_22_port);
   registers_reg_22_21_inst : DLH_X1 port map( G => n2032, D => n2088, Q => 
                           registers_22_21_port);
   registers_reg_22_20_inst : DLH_X1 port map( G => n2031, D => n2091, Q => 
                           registers_22_20_port);
   registers_reg_22_19_inst : DLH_X1 port map( G => n2032, D => n2094, Q => 
                           registers_22_19_port);
   registers_reg_22_18_inst : DLH_X1 port map( G => n2032, D => n2097, Q => 
                           registers_22_18_port);
   registers_reg_22_17_inst : DLH_X1 port map( G => n2031, D => n2100, Q => 
                           registers_22_17_port);
   registers_reg_22_16_inst : DLH_X1 port map( G => n2032, D => n2103, Q => 
                           registers_22_16_port);
   registers_reg_22_15_inst : DLH_X1 port map( G => n2032, D => n2106, Q => 
                           registers_22_15_port);
   registers_reg_22_14_inst : DLH_X1 port map( G => n2032, D => n2109, Q => 
                           registers_22_14_port);
   registers_reg_22_13_inst : DLH_X1 port map( G => n2032, D => n2112, Q => 
                           registers_22_13_port);
   registers_reg_22_12_inst : DLH_X1 port map( G => n2032, D => n2115, Q => 
                           registers_22_12_port);
   registers_reg_22_11_inst : DLH_X1 port map( G => n2033, D => n2118, Q => 
                           registers_22_11_port);
   registers_reg_22_10_inst : DLH_X1 port map( G => n2033, D => n2121, Q => 
                           registers_22_10_port);
   registers_reg_22_9_inst : DLH_X1 port map( G => n2033, D => n2124, Q => 
                           registers_22_9_port);
   registers_reg_22_8_inst : DLH_X1 port map( G => n2033, D => n2127, Q => 
                           registers_22_8_port);
   registers_reg_22_7_inst : DLH_X1 port map( G => n2033, D => n2130, Q => 
                           registers_22_7_port);
   registers_reg_22_6_inst : DLH_X1 port map( G => n2033, D => n2133, Q => 
                           registers_22_6_port);
   registers_reg_22_5_inst : DLH_X1 port map( G => n2033, D => n2136, Q => 
                           registers_22_5_port);
   registers_reg_22_4_inst : DLH_X1 port map( G => n2033, D => n2139, Q => 
                           registers_22_4_port);
   registers_reg_22_3_inst : DLH_X1 port map( G => n2033, D => n2142, Q => 
                           registers_22_3_port);
   registers_reg_22_2_inst : DLH_X1 port map( G => n2033, D => n2145, Q => 
                           registers_22_2_port);
   registers_reg_22_1_inst : DLH_X1 port map( G => n2031, D => n2148, Q => 
                           registers_22_1_port);
   registers_reg_22_0_inst : DLH_X1 port map( G => n2031, D => n2151, Q => 
                           registers_22_0_port);
   registers_reg_23_31_inst : DLH_X1 port map( G => n2034, D => n2058, Q => 
                           registers_23_31_port);
   registers_reg_23_30_inst : DLH_X1 port map( G => n2034, D => n2061, Q => 
                           registers_23_30_port);
   registers_reg_23_29_inst : DLH_X1 port map( G => n2034, D => n2064, Q => 
                           registers_23_29_port);
   registers_reg_23_28_inst : DLH_X1 port map( G => n2034, D => n2067, Q => 
                           registers_23_28_port);
   registers_reg_23_27_inst : DLH_X1 port map( G => n2034, D => n2070, Q => 
                           registers_23_27_port);
   registers_reg_23_26_inst : DLH_X1 port map( G => n2034, D => n2073, Q => 
                           registers_23_26_port);
   registers_reg_23_25_inst : DLH_X1 port map( G => n2034, D => n2076, Q => 
                           registers_23_25_port);
   registers_reg_23_24_inst : DLH_X1 port map( G => n2035, D => n2079, Q => 
                           registers_23_24_port);
   registers_reg_23_23_inst : DLH_X1 port map( G => n2035, D => n2082, Q => 
                           registers_23_23_port);
   registers_reg_23_22_inst : DLH_X1 port map( G => n2035, D => n2085, Q => 
                           registers_23_22_port);
   registers_reg_23_21_inst : DLH_X1 port map( G => n2035, D => n2088, Q => 
                           registers_23_21_port);
   registers_reg_23_20_inst : DLH_X1 port map( G => n2034, D => n2091, Q => 
                           registers_23_20_port);
   registers_reg_23_19_inst : DLH_X1 port map( G => n2035, D => n2094, Q => 
                           registers_23_19_port);
   registers_reg_23_18_inst : DLH_X1 port map( G => n2035, D => n2097, Q => 
                           registers_23_18_port);
   registers_reg_23_17_inst : DLH_X1 port map( G => n2034, D => n2100, Q => 
                           registers_23_17_port);
   registers_reg_23_16_inst : DLH_X1 port map( G => n2035, D => n2103, Q => 
                           registers_23_16_port);
   registers_reg_23_15_inst : DLH_X1 port map( G => n2035, D => n2106, Q => 
                           registers_23_15_port);
   registers_reg_23_14_inst : DLH_X1 port map( G => n2035, D => n2109, Q => 
                           registers_23_14_port);
   registers_reg_23_13_inst : DLH_X1 port map( G => n2035, D => n2112, Q => 
                           registers_23_13_port);
   registers_reg_23_12_inst : DLH_X1 port map( G => n2035, D => n2115, Q => 
                           registers_23_12_port);
   registers_reg_23_11_inst : DLH_X1 port map( G => n2036, D => n2118, Q => 
                           registers_23_11_port);
   registers_reg_23_10_inst : DLH_X1 port map( G => n2036, D => n2121, Q => 
                           registers_23_10_port);
   registers_reg_23_9_inst : DLH_X1 port map( G => n2036, D => n2124, Q => 
                           registers_23_9_port);
   registers_reg_23_8_inst : DLH_X1 port map( G => n2036, D => n2127, Q => 
                           registers_23_8_port);
   registers_reg_23_7_inst : DLH_X1 port map( G => n2036, D => n2130, Q => 
                           registers_23_7_port);
   registers_reg_23_6_inst : DLH_X1 port map( G => n2036, D => n2133, Q => 
                           registers_23_6_port);
   registers_reg_23_5_inst : DLH_X1 port map( G => n2036, D => n2136, Q => 
                           registers_23_5_port);
   registers_reg_23_4_inst : DLH_X1 port map( G => n2036, D => n2139, Q => 
                           registers_23_4_port);
   registers_reg_23_3_inst : DLH_X1 port map( G => n2036, D => n2142, Q => 
                           registers_23_3_port);
   registers_reg_23_2_inst : DLH_X1 port map( G => n2036, D => n2145, Q => 
                           registers_23_2_port);
   registers_reg_23_1_inst : DLH_X1 port map( G => n2034, D => n2148, Q => 
                           registers_23_1_port);
   registers_reg_23_0_inst : DLH_X1 port map( G => n2034, D => n2151, Q => 
                           registers_23_0_port);
   registers_reg_24_31_inst : DLH_X1 port map( G => n2037, D => n2058, Q => 
                           registers_24_31_port);
   registers_reg_24_30_inst : DLH_X1 port map( G => n2037, D => n2061, Q => 
                           registers_24_30_port);
   registers_reg_24_29_inst : DLH_X1 port map( G => n2037, D => n2064, Q => 
                           registers_24_29_port);
   registers_reg_24_28_inst : DLH_X1 port map( G => n2037, D => n2067, Q => 
                           registers_24_28_port);
   registers_reg_24_27_inst : DLH_X1 port map( G => n2037, D => n2070, Q => 
                           registers_24_27_port);
   registers_reg_24_26_inst : DLH_X1 port map( G => n2037, D => n2073, Q => 
                           registers_24_26_port);
   registers_reg_24_25_inst : DLH_X1 port map( G => n2037, D => n2076, Q => 
                           registers_24_25_port);
   registers_reg_24_24_inst : DLH_X1 port map( G => n2038, D => n2079, Q => 
                           registers_24_24_port);
   registers_reg_24_23_inst : DLH_X1 port map( G => n2038, D => n2082, Q => 
                           registers_24_23_port);
   registers_reg_24_22_inst : DLH_X1 port map( G => n2038, D => n2085, Q => 
                           registers_24_22_port);
   registers_reg_24_21_inst : DLH_X1 port map( G => n2038, D => n2088, Q => 
                           registers_24_21_port);
   registers_reg_24_20_inst : DLH_X1 port map( G => n2037, D => n2091, Q => 
                           registers_24_20_port);
   registers_reg_24_19_inst : DLH_X1 port map( G => n2038, D => n2094, Q => 
                           registers_24_19_port);
   registers_reg_24_18_inst : DLH_X1 port map( G => n2038, D => n2097, Q => 
                           registers_24_18_port);
   registers_reg_24_17_inst : DLH_X1 port map( G => n2037, D => n2100, Q => 
                           registers_24_17_port);
   registers_reg_24_16_inst : DLH_X1 port map( G => n2038, D => n2103, Q => 
                           registers_24_16_port);
   registers_reg_24_15_inst : DLH_X1 port map( G => n2038, D => n2106, Q => 
                           registers_24_15_port);
   registers_reg_24_14_inst : DLH_X1 port map( G => n2038, D => n2109, Q => 
                           registers_24_14_port);
   registers_reg_24_13_inst : DLH_X1 port map( G => n2038, D => n2112, Q => 
                           registers_24_13_port);
   registers_reg_24_12_inst : DLH_X1 port map( G => n2038, D => n2115, Q => 
                           registers_24_12_port);
   registers_reg_24_11_inst : DLH_X1 port map( G => n2039, D => n2118, Q => 
                           registers_24_11_port);
   registers_reg_24_10_inst : DLH_X1 port map( G => n2039, D => n2121, Q => 
                           registers_24_10_port);
   registers_reg_24_9_inst : DLH_X1 port map( G => n2039, D => n2124, Q => 
                           registers_24_9_port);
   registers_reg_24_8_inst : DLH_X1 port map( G => n2039, D => n2127, Q => 
                           registers_24_8_port);
   registers_reg_24_7_inst : DLH_X1 port map( G => n2039, D => n2130, Q => 
                           registers_24_7_port);
   registers_reg_24_6_inst : DLH_X1 port map( G => n2039, D => n2133, Q => 
                           registers_24_6_port);
   registers_reg_24_5_inst : DLH_X1 port map( G => n2039, D => n2136, Q => 
                           registers_24_5_port);
   registers_reg_24_4_inst : DLH_X1 port map( G => n2039, D => n2139, Q => 
                           registers_24_4_port);
   registers_reg_24_3_inst : DLH_X1 port map( G => n2039, D => n2142, Q => 
                           registers_24_3_port);
   registers_reg_24_2_inst : DLH_X1 port map( G => n2039, D => n2145, Q => 
                           registers_24_2_port);
   registers_reg_24_1_inst : DLH_X1 port map( G => n2037, D => n2148, Q => 
                           registers_24_1_port);
   registers_reg_24_0_inst : DLH_X1 port map( G => n2037, D => n2151, Q => 
                           registers_24_0_port);
   registers_reg_25_31_inst : DLH_X1 port map( G => n2040, D => n2058, Q => 
                           registers_25_31_port);
   registers_reg_25_30_inst : DLH_X1 port map( G => n2040, D => n2061, Q => 
                           registers_25_30_port);
   registers_reg_25_29_inst : DLH_X1 port map( G => n2040, D => n2064, Q => 
                           registers_25_29_port);
   registers_reg_25_28_inst : DLH_X1 port map( G => n2040, D => n2067, Q => 
                           registers_25_28_port);
   registers_reg_25_27_inst : DLH_X1 port map( G => n2040, D => n2070, Q => 
                           registers_25_27_port);
   registers_reg_25_26_inst : DLH_X1 port map( G => n2040, D => n2073, Q => 
                           registers_25_26_port);
   registers_reg_25_25_inst : DLH_X1 port map( G => n2040, D => n2076, Q => 
                           registers_25_25_port);
   registers_reg_25_24_inst : DLH_X1 port map( G => n2041, D => n2079, Q => 
                           registers_25_24_port);
   registers_reg_25_23_inst : DLH_X1 port map( G => n2041, D => n2082, Q => 
                           registers_25_23_port);
   registers_reg_25_22_inst : DLH_X1 port map( G => n2041, D => n2085, Q => 
                           registers_25_22_port);
   registers_reg_25_21_inst : DLH_X1 port map( G => n2041, D => n2088, Q => 
                           registers_25_21_port);
   registers_reg_25_20_inst : DLH_X1 port map( G => n2040, D => n2091, Q => 
                           registers_25_20_port);
   registers_reg_25_19_inst : DLH_X1 port map( G => n2041, D => n2094, Q => 
                           registers_25_19_port);
   registers_reg_25_18_inst : DLH_X1 port map( G => n2041, D => n2097, Q => 
                           registers_25_18_port);
   registers_reg_25_17_inst : DLH_X1 port map( G => n2040, D => n2100, Q => 
                           registers_25_17_port);
   registers_reg_25_16_inst : DLH_X1 port map( G => n2041, D => n2103, Q => 
                           registers_25_16_port);
   registers_reg_25_15_inst : DLH_X1 port map( G => n2041, D => n2106, Q => 
                           registers_25_15_port);
   registers_reg_25_14_inst : DLH_X1 port map( G => n2041, D => n2109, Q => 
                           registers_25_14_port);
   registers_reg_25_13_inst : DLH_X1 port map( G => n2041, D => n2112, Q => 
                           registers_25_13_port);
   registers_reg_25_12_inst : DLH_X1 port map( G => n2041, D => n2115, Q => 
                           registers_25_12_port);
   registers_reg_25_11_inst : DLH_X1 port map( G => n2042, D => n2118, Q => 
                           registers_25_11_port);
   registers_reg_25_10_inst : DLH_X1 port map( G => n2042, D => n2121, Q => 
                           registers_25_10_port);
   registers_reg_25_9_inst : DLH_X1 port map( G => n2042, D => n2124, Q => 
                           registers_25_9_port);
   registers_reg_25_8_inst : DLH_X1 port map( G => n2042, D => n2127, Q => 
                           registers_25_8_port);
   registers_reg_25_7_inst : DLH_X1 port map( G => n2042, D => n2130, Q => 
                           registers_25_7_port);
   registers_reg_25_6_inst : DLH_X1 port map( G => n2042, D => n2133, Q => 
                           registers_25_6_port);
   registers_reg_25_5_inst : DLH_X1 port map( G => n2042, D => n2136, Q => 
                           registers_25_5_port);
   registers_reg_25_4_inst : DLH_X1 port map( G => n2042, D => n2139, Q => 
                           registers_25_4_port);
   registers_reg_25_3_inst : DLH_X1 port map( G => n2042, D => n2142, Q => 
                           registers_25_3_port);
   registers_reg_25_2_inst : DLH_X1 port map( G => n2042, D => n2145, Q => 
                           registers_25_2_port);
   registers_reg_25_1_inst : DLH_X1 port map( G => n2040, D => n2148, Q => 
                           registers_25_1_port);
   registers_reg_25_0_inst : DLH_X1 port map( G => n2040, D => n2151, Q => 
                           registers_25_0_port);
   registers_reg_26_31_inst : DLH_X1 port map( G => n2043, D => n2058, Q => 
                           registers_26_31_port);
   registers_reg_26_30_inst : DLH_X1 port map( G => n2043, D => n2061, Q => 
                           registers_26_30_port);
   registers_reg_26_29_inst : DLH_X1 port map( G => n2043, D => n2064, Q => 
                           registers_26_29_port);
   registers_reg_26_28_inst : DLH_X1 port map( G => n2043, D => n2067, Q => 
                           registers_26_28_port);
   registers_reg_26_27_inst : DLH_X1 port map( G => n2043, D => n2070, Q => 
                           registers_26_27_port);
   registers_reg_26_26_inst : DLH_X1 port map( G => n2043, D => n2073, Q => 
                           registers_26_26_port);
   registers_reg_26_25_inst : DLH_X1 port map( G => n2043, D => n2076, Q => 
                           registers_26_25_port);
   registers_reg_26_24_inst : DLH_X1 port map( G => n2044, D => n2079, Q => 
                           registers_26_24_port);
   registers_reg_26_23_inst : DLH_X1 port map( G => n2044, D => n2082, Q => 
                           registers_26_23_port);
   registers_reg_26_22_inst : DLH_X1 port map( G => n2044, D => n2085, Q => 
                           registers_26_22_port);
   registers_reg_26_21_inst : DLH_X1 port map( G => n2044, D => n2088, Q => 
                           registers_26_21_port);
   registers_reg_26_20_inst : DLH_X1 port map( G => n2043, D => n2091, Q => 
                           registers_26_20_port);
   registers_reg_26_19_inst : DLH_X1 port map( G => n2044, D => n2094, Q => 
                           registers_26_19_port);
   registers_reg_26_18_inst : DLH_X1 port map( G => n2044, D => n2097, Q => 
                           registers_26_18_port);
   registers_reg_26_17_inst : DLH_X1 port map( G => n2043, D => n2100, Q => 
                           registers_26_17_port);
   registers_reg_26_16_inst : DLH_X1 port map( G => n2044, D => n2103, Q => 
                           registers_26_16_port);
   registers_reg_26_15_inst : DLH_X1 port map( G => n2044, D => n2106, Q => 
                           registers_26_15_port);
   registers_reg_26_14_inst : DLH_X1 port map( G => n2044, D => n2109, Q => 
                           registers_26_14_port);
   registers_reg_26_13_inst : DLH_X1 port map( G => n2044, D => n2112, Q => 
                           registers_26_13_port);
   registers_reg_26_12_inst : DLH_X1 port map( G => n2044, D => n2115, Q => 
                           registers_26_12_port);
   registers_reg_26_11_inst : DLH_X1 port map( G => n2045, D => n2118, Q => 
                           registers_26_11_port);
   registers_reg_26_10_inst : DLH_X1 port map( G => n2045, D => n2121, Q => 
                           registers_26_10_port);
   registers_reg_26_9_inst : DLH_X1 port map( G => n2045, D => n2124, Q => 
                           registers_26_9_port);
   registers_reg_26_8_inst : DLH_X1 port map( G => n2045, D => n2127, Q => 
                           registers_26_8_port);
   registers_reg_26_7_inst : DLH_X1 port map( G => n2045, D => n2130, Q => 
                           registers_26_7_port);
   registers_reg_26_6_inst : DLH_X1 port map( G => n2045, D => n2133, Q => 
                           registers_26_6_port);
   registers_reg_26_5_inst : DLH_X1 port map( G => n2045, D => n2136, Q => 
                           registers_26_5_port);
   registers_reg_26_4_inst : DLH_X1 port map( G => n2045, D => n2139, Q => 
                           registers_26_4_port);
   registers_reg_26_3_inst : DLH_X1 port map( G => n2045, D => n2142, Q => 
                           registers_26_3_port);
   registers_reg_26_2_inst : DLH_X1 port map( G => n2045, D => n2145, Q => 
                           registers_26_2_port);
   registers_reg_26_1_inst : DLH_X1 port map( G => n2043, D => n2148, Q => 
                           registers_26_1_port);
   registers_reg_26_0_inst : DLH_X1 port map( G => n2043, D => n2151, Q => 
                           registers_26_0_port);
   registers_reg_27_31_inst : DLH_X1 port map( G => n2046, D => n2058, Q => 
                           registers_27_31_port);
   registers_reg_27_30_inst : DLH_X1 port map( G => n2046, D => n2061, Q => 
                           registers_27_30_port);
   registers_reg_27_29_inst : DLH_X1 port map( G => n2046, D => n2064, Q => 
                           registers_27_29_port);
   registers_reg_27_28_inst : DLH_X1 port map( G => n2046, D => n2067, Q => 
                           registers_27_28_port);
   registers_reg_27_27_inst : DLH_X1 port map( G => n2046, D => n2070, Q => 
                           registers_27_27_port);
   registers_reg_27_26_inst : DLH_X1 port map( G => n2046, D => n2073, Q => 
                           registers_27_26_port);
   registers_reg_27_25_inst : DLH_X1 port map( G => n2046, D => n2076, Q => 
                           registers_27_25_port);
   registers_reg_27_24_inst : DLH_X1 port map( G => n2047, D => n2079, Q => 
                           registers_27_24_port);
   registers_reg_27_23_inst : DLH_X1 port map( G => n2047, D => n2082, Q => 
                           registers_27_23_port);
   registers_reg_27_22_inst : DLH_X1 port map( G => n2047, D => n2085, Q => 
                           registers_27_22_port);
   registers_reg_27_21_inst : DLH_X1 port map( G => n2047, D => n2088, Q => 
                           registers_27_21_port);
   registers_reg_27_20_inst : DLH_X1 port map( G => n2046, D => n2091, Q => 
                           registers_27_20_port);
   registers_reg_27_19_inst : DLH_X1 port map( G => n2047, D => n2094, Q => 
                           registers_27_19_port);
   registers_reg_27_18_inst : DLH_X1 port map( G => n2047, D => n2097, Q => 
                           registers_27_18_port);
   registers_reg_27_17_inst : DLH_X1 port map( G => n2046, D => n2100, Q => 
                           registers_27_17_port);
   registers_reg_27_16_inst : DLH_X1 port map( G => n2047, D => n2103, Q => 
                           registers_27_16_port);
   registers_reg_27_15_inst : DLH_X1 port map( G => n2047, D => n2106, Q => 
                           registers_27_15_port);
   registers_reg_27_14_inst : DLH_X1 port map( G => n2047, D => n2109, Q => 
                           registers_27_14_port);
   registers_reg_27_13_inst : DLH_X1 port map( G => n2047, D => n2112, Q => 
                           registers_27_13_port);
   registers_reg_27_12_inst : DLH_X1 port map( G => n2047, D => n2115, Q => 
                           registers_27_12_port);
   registers_reg_27_11_inst : DLH_X1 port map( G => n2048, D => n2118, Q => 
                           registers_27_11_port);
   registers_reg_27_10_inst : DLH_X1 port map( G => n2048, D => n2121, Q => 
                           registers_27_10_port);
   registers_reg_27_9_inst : DLH_X1 port map( G => n2048, D => n2124, Q => 
                           registers_27_9_port);
   registers_reg_27_8_inst : DLH_X1 port map( G => n2048, D => n2127, Q => 
                           registers_27_8_port);
   registers_reg_27_7_inst : DLH_X1 port map( G => n2048, D => n2130, Q => 
                           registers_27_7_port);
   registers_reg_27_6_inst : DLH_X1 port map( G => n2048, D => n2133, Q => 
                           registers_27_6_port);
   registers_reg_27_5_inst : DLH_X1 port map( G => n2048, D => n2136, Q => 
                           registers_27_5_port);
   registers_reg_27_4_inst : DLH_X1 port map( G => n2048, D => n2139, Q => 
                           registers_27_4_port);
   registers_reg_27_3_inst : DLH_X1 port map( G => n2048, D => n2142, Q => 
                           registers_27_3_port);
   registers_reg_27_2_inst : DLH_X1 port map( G => n2048, D => n2145, Q => 
                           registers_27_2_port);
   registers_reg_27_1_inst : DLH_X1 port map( G => n2046, D => n2148, Q => 
                           registers_27_1_port);
   registers_reg_27_0_inst : DLH_X1 port map( G => n2046, D => n2151, Q => 
                           registers_27_0_port);
   registers_reg_28_31_inst : DLH_X1 port map( G => n2049, D => n2058, Q => 
                           registers_28_31_port);
   registers_reg_28_30_inst : DLH_X1 port map( G => n2049, D => n2061, Q => 
                           registers_28_30_port);
   registers_reg_28_29_inst : DLH_X1 port map( G => n2049, D => n2064, Q => 
                           registers_28_29_port);
   registers_reg_28_28_inst : DLH_X1 port map( G => n2049, D => n2067, Q => 
                           registers_28_28_port);
   registers_reg_28_27_inst : DLH_X1 port map( G => n2049, D => n2070, Q => 
                           registers_28_27_port);
   registers_reg_28_26_inst : DLH_X1 port map( G => n2049, D => n2073, Q => 
                           registers_28_26_port);
   registers_reg_28_25_inst : DLH_X1 port map( G => n2049, D => n2076, Q => 
                           registers_28_25_port);
   registers_reg_28_24_inst : DLH_X1 port map( G => n2050, D => n2079, Q => 
                           registers_28_24_port);
   registers_reg_28_23_inst : DLH_X1 port map( G => n2050, D => n2082, Q => 
                           registers_28_23_port);
   registers_reg_28_22_inst : DLH_X1 port map( G => n2050, D => n2085, Q => 
                           registers_28_22_port);
   registers_reg_28_21_inst : DLH_X1 port map( G => n2050, D => n2088, Q => 
                           registers_28_21_port);
   registers_reg_28_20_inst : DLH_X1 port map( G => n2049, D => n2091, Q => 
                           registers_28_20_port);
   registers_reg_28_19_inst : DLH_X1 port map( G => n2050, D => n2094, Q => 
                           registers_28_19_port);
   registers_reg_28_18_inst : DLH_X1 port map( G => n2050, D => n2097, Q => 
                           registers_28_18_port);
   registers_reg_28_17_inst : DLH_X1 port map( G => n2049, D => n2100, Q => 
                           registers_28_17_port);
   registers_reg_28_16_inst : DLH_X1 port map( G => n2050, D => n2103, Q => 
                           registers_28_16_port);
   registers_reg_28_15_inst : DLH_X1 port map( G => n2050, D => n2106, Q => 
                           registers_28_15_port);
   registers_reg_28_14_inst : DLH_X1 port map( G => n2050, D => n2109, Q => 
                           registers_28_14_port);
   registers_reg_28_13_inst : DLH_X1 port map( G => n2050, D => n2112, Q => 
                           registers_28_13_port);
   registers_reg_28_12_inst : DLH_X1 port map( G => n2050, D => n2115, Q => 
                           registers_28_12_port);
   registers_reg_28_11_inst : DLH_X1 port map( G => n2051, D => n2118, Q => 
                           registers_28_11_port);
   registers_reg_28_10_inst : DLH_X1 port map( G => n2051, D => n2121, Q => 
                           registers_28_10_port);
   registers_reg_28_9_inst : DLH_X1 port map( G => n2051, D => n2124, Q => 
                           registers_28_9_port);
   registers_reg_28_8_inst : DLH_X1 port map( G => n2051, D => n2127, Q => 
                           registers_28_8_port);
   registers_reg_28_7_inst : DLH_X1 port map( G => n2051, D => n2130, Q => 
                           registers_28_7_port);
   registers_reg_28_6_inst : DLH_X1 port map( G => n2051, D => n2133, Q => 
                           registers_28_6_port);
   registers_reg_28_5_inst : DLH_X1 port map( G => n2051, D => n2136, Q => 
                           registers_28_5_port);
   registers_reg_28_4_inst : DLH_X1 port map( G => n2051, D => n2139, Q => 
                           registers_28_4_port);
   registers_reg_28_3_inst : DLH_X1 port map( G => n2051, D => n2142, Q => 
                           registers_28_3_port);
   registers_reg_28_2_inst : DLH_X1 port map( G => n2051, D => n2145, Q => 
                           registers_28_2_port);
   registers_reg_28_1_inst : DLH_X1 port map( G => n2049, D => n2148, Q => 
                           registers_28_1_port);
   registers_reg_28_0_inst : DLH_X1 port map( G => n2049, D => n2151, Q => 
                           registers_28_0_port);
   registers_reg_29_31_inst : DLH_X1 port map( G => n2052, D => n2058, Q => 
                           registers_29_31_port);
   registers_reg_29_30_inst : DLH_X1 port map( G => n2052, D => n2061, Q => 
                           registers_29_30_port);
   registers_reg_29_29_inst : DLH_X1 port map( G => n2052, D => n2064, Q => 
                           registers_29_29_port);
   registers_reg_29_28_inst : DLH_X1 port map( G => n2052, D => n2067, Q => 
                           registers_29_28_port);
   registers_reg_29_27_inst : DLH_X1 port map( G => n2052, D => n2070, Q => 
                           registers_29_27_port);
   registers_reg_29_26_inst : DLH_X1 port map( G => n2052, D => n2073, Q => 
                           registers_29_26_port);
   registers_reg_29_25_inst : DLH_X1 port map( G => n2052, D => n2076, Q => 
                           registers_29_25_port);
   registers_reg_29_24_inst : DLH_X1 port map( G => n2053, D => n2079, Q => 
                           registers_29_24_port);
   registers_reg_29_23_inst : DLH_X1 port map( G => n2053, D => n2082, Q => 
                           registers_29_23_port);
   registers_reg_29_22_inst : DLH_X1 port map( G => n2053, D => n2085, Q => 
                           registers_29_22_port);
   registers_reg_29_21_inst : DLH_X1 port map( G => n2053, D => n2088, Q => 
                           registers_29_21_port);
   registers_reg_29_20_inst : DLH_X1 port map( G => n2052, D => n2091, Q => 
                           registers_29_20_port);
   registers_reg_29_19_inst : DLH_X1 port map( G => n2053, D => n2094, Q => 
                           registers_29_19_port);
   registers_reg_29_18_inst : DLH_X1 port map( G => n2053, D => n2097, Q => 
                           registers_29_18_port);
   registers_reg_29_17_inst : DLH_X1 port map( G => n2052, D => n2100, Q => 
                           registers_29_17_port);
   registers_reg_29_16_inst : DLH_X1 port map( G => n2053, D => n2103, Q => 
                           registers_29_16_port);
   registers_reg_29_15_inst : DLH_X1 port map( G => n2053, D => n2106, Q => 
                           registers_29_15_port);
   registers_reg_29_14_inst : DLH_X1 port map( G => n2053, D => n2109, Q => 
                           registers_29_14_port);
   registers_reg_29_13_inst : DLH_X1 port map( G => n2053, D => n2112, Q => 
                           registers_29_13_port);
   registers_reg_29_12_inst : DLH_X1 port map( G => n2053, D => n2115, Q => 
                           registers_29_12_port);
   registers_reg_29_11_inst : DLH_X1 port map( G => n2054, D => n2118, Q => 
                           registers_29_11_port);
   registers_reg_29_10_inst : DLH_X1 port map( G => n2054, D => n2121, Q => 
                           registers_29_10_port);
   registers_reg_29_9_inst : DLH_X1 port map( G => n2054, D => n2124, Q => 
                           registers_29_9_port);
   registers_reg_29_8_inst : DLH_X1 port map( G => n2054, D => n2127, Q => 
                           registers_29_8_port);
   registers_reg_29_7_inst : DLH_X1 port map( G => n2054, D => n2130, Q => 
                           registers_29_7_port);
   registers_reg_29_6_inst : DLH_X1 port map( G => n2054, D => n2133, Q => 
                           registers_29_6_port);
   registers_reg_29_5_inst : DLH_X1 port map( G => n2054, D => n2136, Q => 
                           registers_29_5_port);
   registers_reg_29_4_inst : DLH_X1 port map( G => n2054, D => n2139, Q => 
                           registers_29_4_port);
   registers_reg_29_3_inst : DLH_X1 port map( G => n2054, D => n2142, Q => 
                           registers_29_3_port);
   registers_reg_29_2_inst : DLH_X1 port map( G => n2054, D => n2145, Q => 
                           registers_29_2_port);
   registers_reg_29_1_inst : DLH_X1 port map( G => n2052, D => n2148, Q => 
                           registers_29_1_port);
   registers_reg_29_0_inst : DLH_X1 port map( G => n2052, D => n2151, Q => 
                           registers_29_0_port);
   registers_reg_30_31_inst : DLH_X1 port map( G => n2055, D => n2058, Q => 
                           registers_30_31_port);
   registers_reg_30_30_inst : DLH_X1 port map( G => n2055, D => n2061, Q => 
                           registers_30_30_port);
   registers_reg_30_29_inst : DLH_X1 port map( G => n2055, D => n2064, Q => 
                           registers_30_29_port);
   registers_reg_30_28_inst : DLH_X1 port map( G => n2055, D => n2067, Q => 
                           registers_30_28_port);
   registers_reg_30_27_inst : DLH_X1 port map( G => n2055, D => n2070, Q => 
                           registers_30_27_port);
   registers_reg_30_26_inst : DLH_X1 port map( G => n2055, D => n2073, Q => 
                           registers_30_26_port);
   registers_reg_30_25_inst : DLH_X1 port map( G => n2055, D => n2076, Q => 
                           registers_30_25_port);
   registers_reg_30_24_inst : DLH_X1 port map( G => n2056, D => n2079, Q => 
                           registers_30_24_port);
   registers_reg_30_23_inst : DLH_X1 port map( G => n2056, D => n2082, Q => 
                           registers_30_23_port);
   registers_reg_30_22_inst : DLH_X1 port map( G => n2056, D => n2085, Q => 
                           registers_30_22_port);
   registers_reg_30_21_inst : DLH_X1 port map( G => n2056, D => n2088, Q => 
                           registers_30_21_port);
   registers_reg_30_20_inst : DLH_X1 port map( G => n2055, D => n2091, Q => 
                           registers_30_20_port);
   registers_reg_30_19_inst : DLH_X1 port map( G => n2056, D => n2094, Q => 
                           registers_30_19_port);
   registers_reg_30_18_inst : DLH_X1 port map( G => n2056, D => n2097, Q => 
                           registers_30_18_port);
   registers_reg_30_17_inst : DLH_X1 port map( G => n2055, D => n2100, Q => 
                           registers_30_17_port);
   registers_reg_30_16_inst : DLH_X1 port map( G => n2056, D => n2103, Q => 
                           registers_30_16_port);
   registers_reg_30_15_inst : DLH_X1 port map( G => n2056, D => n2106, Q => 
                           registers_30_15_port);
   registers_reg_30_14_inst : DLH_X1 port map( G => n2056, D => n2109, Q => 
                           registers_30_14_port);
   registers_reg_30_13_inst : DLH_X1 port map( G => n2056, D => n2112, Q => 
                           registers_30_13_port);
   registers_reg_30_12_inst : DLH_X1 port map( G => n2056, D => n2115, Q => 
                           registers_30_12_port);
   registers_reg_30_11_inst : DLH_X1 port map( G => n2057, D => n2118, Q => 
                           registers_30_11_port);
   registers_reg_30_10_inst : DLH_X1 port map( G => n2057, D => n2121, Q => 
                           registers_30_10_port);
   registers_reg_30_9_inst : DLH_X1 port map( G => n2057, D => n2124, Q => 
                           registers_30_9_port);
   registers_reg_30_8_inst : DLH_X1 port map( G => n2057, D => n2127, Q => 
                           registers_30_8_port);
   registers_reg_30_7_inst : DLH_X1 port map( G => n2057, D => n2130, Q => 
                           registers_30_7_port);
   registers_reg_30_6_inst : DLH_X1 port map( G => n2057, D => n2133, Q => 
                           registers_30_6_port);
   registers_reg_30_5_inst : DLH_X1 port map( G => n2057, D => n2136, Q => 
                           registers_30_5_port);
   registers_reg_30_4_inst : DLH_X1 port map( G => n2057, D => n2139, Q => 
                           registers_30_4_port);
   registers_reg_30_3_inst : DLH_X1 port map( G => n2057, D => n2142, Q => 
                           registers_30_3_port);
   registers_reg_30_2_inst : DLH_X1 port map( G => n2057, D => n2145, Q => 
                           registers_30_2_port);
   registers_reg_30_1_inst : DLH_X1 port map( G => n2055, D => n2148, Q => 
                           registers_30_1_port);
   registers_reg_30_0_inst : DLH_X1 port map( G => n2055, D => n2151, Q => 
                           registers_30_0_port);
   registers_reg_31_31_inst : DLH_X1 port map( G => n2154, D => n2058, Q => 
                           registers_31_31_port);
   registers_reg_31_30_inst : DLH_X1 port map( G => n2154, D => n2061, Q => 
                           registers_31_30_port);
   registers_reg_31_29_inst : DLH_X1 port map( G => n2154, D => n2064, Q => 
                           registers_31_29_port);
   registers_reg_31_28_inst : DLH_X1 port map( G => n2154, D => n2067, Q => 
                           registers_31_28_port);
   registers_reg_31_27_inst : DLH_X1 port map( G => n2154, D => n2070, Q => 
                           registers_31_27_port);
   registers_reg_31_26_inst : DLH_X1 port map( G => n2154, D => n2073, Q => 
                           registers_31_26_port);
   registers_reg_31_25_inst : DLH_X1 port map( G => n2154, D => n2076, Q => 
                           registers_31_25_port);
   registers_reg_31_24_inst : DLH_X1 port map( G => n2155, D => n2079, Q => 
                           registers_31_24_port);
   registers_reg_31_23_inst : DLH_X1 port map( G => n2155, D => n2082, Q => 
                           registers_31_23_port);
   registers_reg_31_22_inst : DLH_X1 port map( G => n2155, D => n2085, Q => 
                           registers_31_22_port);
   registers_reg_31_21_inst : DLH_X1 port map( G => n2155, D => n2088, Q => 
                           registers_31_21_port);
   registers_reg_31_20_inst : DLH_X1 port map( G => n2154, D => n2091, Q => 
                           registers_31_20_port);
   registers_reg_31_19_inst : DLH_X1 port map( G => n2155, D => n2094, Q => 
                           registers_31_19_port);
   registers_reg_31_18_inst : DLH_X1 port map( G => n2155, D => n2097, Q => 
                           registers_31_18_port);
   registers_reg_31_17_inst : DLH_X1 port map( G => n2154, D => n2100, Q => 
                           registers_31_17_port);
   registers_reg_31_16_inst : DLH_X1 port map( G => n2155, D => n2103, Q => 
                           registers_31_16_port);
   registers_reg_31_15_inst : DLH_X1 port map( G => n2155, D => n2106, Q => 
                           registers_31_15_port);
   registers_reg_31_14_inst : DLH_X1 port map( G => n2155, D => n2109, Q => 
                           registers_31_14_port);
   registers_reg_31_13_inst : DLH_X1 port map( G => n2155, D => n2112, Q => 
                           registers_31_13_port);
   registers_reg_31_12_inst : DLH_X1 port map( G => n2155, D => n2115, Q => 
                           registers_31_12_port);
   registers_reg_31_11_inst : DLH_X1 port map( G => n2156, D => n2118, Q => 
                           registers_31_11_port);
   registers_reg_31_10_inst : DLH_X1 port map( G => n2156, D => n2121, Q => 
                           registers_31_10_port);
   registers_reg_31_9_inst : DLH_X1 port map( G => n2156, D => n2124, Q => 
                           registers_31_9_port);
   registers_reg_31_8_inst : DLH_X1 port map( G => n2156, D => n2127, Q => 
                           registers_31_8_port);
   registers_reg_31_7_inst : DLH_X1 port map( G => n2156, D => n2130, Q => 
                           registers_31_7_port);
   registers_reg_31_6_inst : DLH_X1 port map( G => n2156, D => n2133, Q => 
                           registers_31_6_port);
   registers_reg_31_5_inst : DLH_X1 port map( G => n2156, D => n2136, Q => 
                           registers_31_5_port);
   registers_reg_31_4_inst : DLH_X1 port map( G => n2156, D => n2139, Q => 
                           registers_31_4_port);
   registers_reg_31_3_inst : DLH_X1 port map( G => n2156, D => n2142, Q => 
                           registers_31_3_port);
   registers_reg_31_2_inst : DLH_X1 port map( G => n2156, D => n2145, Q => 
                           registers_31_2_port);
   registers_reg_31_1_inst : DLH_X1 port map( G => n2154, D => n2148, Q => 
                           registers_31_1_port);
   registers_reg_31_0_inst : DLH_X1 port map( G => n2154, D => n2151, Q => 
                           registers_31_0_port);
   out2_reg_31_inst : DLH_X1 port map( G => n1962, D => N243, Q => out2(31));
   out2_reg_30_inst : DLH_X1 port map( G => n1962, D => N244, Q => out2(30));
   out2_reg_29_inst : DLH_X1 port map( G => n1962, D => N245, Q => out2(29));
   out2_reg_28_inst : DLH_X1 port map( G => n1963, D => N246, Q => out2(28));
   out2_reg_27_inst : DLH_X1 port map( G => n1962, D => N247, Q => out2(27));
   out2_reg_26_inst : DLH_X1 port map( G => n1963, D => N248, Q => out2(26));
   out2_reg_25_inst : DLH_X1 port map( G => n1963, D => N249, Q => out2(25));
   out2_reg_24_inst : DLH_X1 port map( G => n1964, D => N250, Q => out2(24));
   out2_reg_23_inst : DLH_X1 port map( G => n1964, D => N251, Q => out2(23));
   out2_reg_22_inst : DLH_X1 port map( G => n1964, D => N252, Q => out2(22));
   out2_reg_21_inst : DLH_X1 port map( G => n1965, D => N253, Q => out2(21));
   out2_reg_20_inst : DLH_X1 port map( G => n1963, D => N254, Q => out2(20));
   out2_reg_19_inst : DLH_X1 port map( G => n1964, D => N255, Q => out2(19));
   out2_reg_18_inst : DLH_X1 port map( G => n1964, D => N256, Q => out2(18));
   out2_reg_17_inst : DLH_X1 port map( G => n1962, D => N257, Q => out2(17));
   out2_reg_16_inst : DLH_X1 port map( G => n1964, D => N258, Q => out2(16));
   out2_reg_15_inst : DLH_X1 port map( G => n1965, D => N259, Q => out2(15));
   out2_reg_14_inst : DLH_X1 port map( G => n1965, D => N260, Q => out2(14));
   out2_reg_13_inst : DLH_X1 port map( G => n1965, D => N261, Q => out2(13));
   out2_reg_12_inst : DLH_X1 port map( G => n1965, D => N262, Q => out2(12));
   out2_reg_11_inst : DLH_X1 port map( G => n1966, D => N263, Q => out2(11));
   out2_reg_10_inst : DLH_X1 port map( G => n1966, D => N264, Q => out2(10));
   out2_reg_9_inst : DLH_X1 port map( G => n1966, D => N265, Q => out2(9));
   out2_reg_8_inst : DLH_X1 port map( G => n1966, D => N266, Q => out2(8));
   out2_reg_7_inst : DLH_X1 port map( G => n1966, D => N267, Q => out2(7));
   out2_reg_6_inst : DLH_X1 port map( G => n1967, D => N268, Q => out2(6));
   out2_reg_5_inst : DLH_X1 port map( G => n1967, D => N269, Q => out2(5));
   out2_reg_4_inst : DLH_X1 port map( G => n1967, D => N270, Q => out2(4));
   out2_reg_3_inst : DLH_X1 port map( G => n1966, D => N271, Q => out2(3));
   out2_reg_2_inst : DLH_X1 port map( G => n1967, D => N272, Q => out2(2));
   out2_reg_1_inst : DLH_X1 port map( G => n1963, D => N273, Q => out2(1));
   out2_reg_0_inst : DLH_X1 port map( G => n1962, D => N274, Q => out2(0));
   out1_reg_31_inst : DLH_X1 port map( G => n1962, D => N146, Q => out1(31));
   out1_reg_30_inst : DLH_X1 port map( G => n1962, D => N147, Q => out1(30));
   out1_reg_29_inst : DLH_X1 port map( G => n1962, D => N148, Q => out1(29));
   out1_reg_28_inst : DLH_X1 port map( G => n1963, D => N149, Q => out1(28));
   out1_reg_27_inst : DLH_X1 port map( G => n1963, D => N150, Q => out1(27));
   out1_reg_26_inst : DLH_X1 port map( G => n1963, D => N151, Q => out1(26));
   out1_reg_25_inst : DLH_X1 port map( G => n1963, D => N152, Q => out1(25));
   out1_reg_24_inst : DLH_X1 port map( G => n1964, D => N153, Q => out1(24));
   out1_reg_23_inst : DLH_X1 port map( G => n1964, D => N154, Q => out1(23));
   out1_reg_22_inst : DLH_X1 port map( G => n1964, D => N155, Q => out1(22));
   out1_reg_21_inst : DLH_X1 port map( G => n1965, D => N156, Q => out1(21));
   out1_reg_20_inst : DLH_X1 port map( G => n1963, D => N157, Q => out1(20));
   out1_reg_19_inst : DLH_X1 port map( G => n1964, D => N158, Q => out1(19));
   out1_reg_18_inst : DLH_X1 port map( G => n1965, D => N159, Q => out1(18));
   out1_reg_17_inst : DLH_X1 port map( G => n1962, D => N160, Q => out1(17));
   out1_reg_16_inst : DLH_X1 port map( G => n1964, D => N161, Q => out1(16));
   out1_reg_15_inst : DLH_X1 port map( G => n1965, D => N162, Q => out1(15));
   out1_reg_14_inst : DLH_X1 port map( G => n1965, D => N163, Q => out1(14));
   out1_reg_13_inst : DLH_X1 port map( G => n1965, D => N164, Q => out1(13));
   out1_reg_12_inst : DLH_X1 port map( G => n1965, D => N165, Q => out1(12));
   out1_reg_11_inst : DLH_X1 port map( G => n1966, D => N166, Q => out1(11));
   out1_reg_10_inst : DLH_X1 port map( G => n1966, D => N167, Q => out1(10));
   out1_reg_9_inst : DLH_X1 port map( G => n1966, D => N168, Q => out1(9));
   out1_reg_8_inst : DLH_X1 port map( G => n1966, D => N169, Q => out1(8));
   out1_reg_7_inst : DLH_X1 port map( G => n1967, D => N170, Q => out1(7));
   out1_reg_6_inst : DLH_X1 port map( G => n1967, D => N171, Q => out1(6));
   out1_reg_5_inst : DLH_X1 port map( G => n1967, D => N172, Q => out1(5));
   out1_reg_4_inst : DLH_X1 port map( G => n1967, D => N173, Q => out1(4));
   out1_reg_3_inst : DLH_X1 port map( G => n1966, D => N174, Q => out1(3));
   out1_reg_2_inst : DLH_X1 port map( G => n1967, D => N175, Q => out1(2));
   out1_reg_1_inst : DLH_X1 port map( G => n1963, D => N176, Q => out1(1));
   out1_reg_0_inst : DLH_X1 port map( G => n1962, D => N177, Q => out1(0));
   U1832 : NAND3_X1 port map( A1 => n2165, A2 => n2164, A3 => n535, ZN => n527)
                           ;
   U1833 : NAND3_X1 port map( A1 => n535, A2 => n2164, A3 => add_wr(3), ZN => 
                           n536);
   U1834 : NAND3_X1 port map( A1 => n535, A2 => n2165, A3 => add_wr(4), ZN => 
                           n538);
   U1835 : NAND3_X1 port map( A1 => n2167, A2 => n2166, A3 => n2168, ZN => n537
                           );
   U1836 : NAND3_X1 port map( A1 => n2167, A2 => n2166, A3 => add_wr(0), ZN => 
                           n528);
   U1837 : NAND3_X1 port map( A1 => n2168, A2 => n2166, A3 => add_wr(1), ZN => 
                           n529);
   U1838 : NAND3_X1 port map( A1 => add_wr(0), A2 => n2166, A3 => add_wr(1), ZN
                           => n530);
   U1839 : NAND3_X1 port map( A1 => n2168, A2 => n2167, A3 => add_wr(2), ZN => 
                           n531);
   U1840 : NAND3_X1 port map( A1 => add_wr(0), A2 => n2167, A3 => add_wr(2), ZN
                           => n532);
   U1841 : NAND3_X1 port map( A1 => add_wr(1), A2 => n2168, A3 => add_wr(2), ZN
                           => n533);
   U1842 : NAND3_X1 port map( A1 => add_wr(3), A2 => n535, A3 => add_wr(4), ZN 
                           => n539);
   U1843 : NAND3_X1 port map( A1 => add_wr(1), A2 => add_wr(0), A3 => add_wr(2)
                           , ZN => n534);
   U3 : NOR2_X1 port map( A1 => n2683, A2 => add_rd1(2), ZN => n1697);
   U4 : NOR2_X1 port map( A1 => n2687, A2 => add_rd2(2), ZN => n1110);
   U5 : BUF_X1 port map( A => n2157, Z => n2161);
   U6 : BUF_X1 port map( A => n2157, Z => n2160);
   U7 : BUF_X1 port map( A => n2157, Z => n2159);
   U8 : BUF_X1 port map( A => n2158, Z => n2162);
   U9 : BUF_X1 port map( A => n2158, Z => n2163);
   U10 : BUF_X1 port map( A => reset, Z => n2157);
   U11 : BUF_X1 port map( A => reset, Z => n2158);
   U12 : BUF_X1 port map( A => n579, Z => n1888);
   U13 : BUF_X1 port map( A => n584, Z => n1876);
   U14 : BUF_X1 port map( A => n579, Z => n1887);
   U15 : BUF_X1 port map( A => n584, Z => n1875);
   U16 : BUF_X1 port map( A => n548, Z => n1960);
   U17 : BUF_X1 port map( A => n553, Z => n1948);
   U18 : BUF_X1 port map( A => n548, Z => n1959);
   U19 : BUF_X1 port map( A => n553, Z => n1947);
   U20 : BUF_X1 port map( A => n551, Z => n1954);
   U21 : BUF_X1 port map( A => n556, Z => n1942);
   U22 : BUF_X1 port map( A => n561, Z => n1930);
   U23 : BUF_X1 port map( A => n566, Z => n1918);
   U24 : BUF_X1 port map( A => n576, Z => n1897);
   U25 : BUF_X1 port map( A => n551, Z => n1953);
   U26 : BUF_X1 port map( A => n556, Z => n1941);
   U27 : BUF_X1 port map( A => n561, Z => n1929);
   U28 : BUF_X1 port map( A => n566, Z => n1917);
   U29 : BUF_X1 port map( A => n576, Z => n1896);
   U30 : BUF_X1 port map( A => n558, Z => n1936);
   U31 : BUF_X1 port map( A => n563, Z => n1924);
   U32 : BUF_X1 port map( A => n573, Z => n1903);
   U33 : BUF_X1 port map( A => n558, Z => n1935);
   U34 : BUF_X1 port map( A => n563, Z => n1923);
   U35 : BUF_X1 port map( A => n573, Z => n1902);
   U36 : BUF_X1 port map( A => n568, Z => n1912);
   U37 : BUF_X1 port map( A => n568, Z => n1911);
   U38 : BUF_X1 port map( A => n552, Z => n1951);
   U39 : BUF_X1 port map( A => n557, Z => n1939);
   U40 : BUF_X1 port map( A => n562, Z => n1927);
   U41 : BUF_X1 port map( A => n567, Z => n1915);
   U42 : BUF_X1 port map( A => n577, Z => n1894);
   U43 : BUF_X1 port map( A => n552, Z => n1950);
   U44 : BUF_X1 port map( A => n557, Z => n1938);
   U45 : BUF_X1 port map( A => n562, Z => n1926);
   U46 : BUF_X1 port map( A => n567, Z => n1914);
   U47 : BUF_X1 port map( A => n577, Z => n1893);
   U48 : BUF_X1 port map( A => n1158, Z => n1816);
   U49 : BUF_X1 port map( A => n1158, Z => n1815);
   U50 : BUF_X1 port map( A => n1168, Z => n1792);
   U51 : BUF_X1 port map( A => n1173, Z => n1780);
   U52 : BUF_X1 port map( A => n1168, Z => n1791);
   U53 : BUF_X1 port map( A => n1173, Z => n1779);
   U54 : BUF_X1 port map( A => n1169, Z => n1789);
   U55 : BUF_X1 port map( A => n1174, Z => n1777);
   U56 : BUF_X1 port map( A => n1169, Z => n1788);
   U57 : BUF_X1 port map( A => n1174, Z => n1776);
   U58 : BUF_X1 port map( A => n1159, Z => n1813);
   U59 : BUF_X1 port map( A => n1159, Z => n1812);
   U60 : BUF_X1 port map( A => n1161, Z => n1807);
   U61 : BUF_X1 port map( A => n1161, Z => n1806);
   U62 : BUF_X1 port map( A => n1136, Z => n1864);
   U63 : BUF_X1 port map( A => n1141, Z => n1852);
   U64 : BUF_X1 port map( A => n1146, Z => n1840);
   U65 : BUF_X1 port map( A => n1151, Z => n1828);
   U66 : BUF_X1 port map( A => n1136, Z => n1863);
   U67 : BUF_X1 port map( A => n1141, Z => n1851);
   U68 : BUF_X1 port map( A => n1146, Z => n1839);
   U69 : BUF_X1 port map( A => n1151, Z => n1827);
   U70 : BUF_X1 port map( A => n1165, Z => n1798);
   U71 : BUF_X1 port map( A => n1170, Z => n1786);
   U72 : BUF_X1 port map( A => n1165, Z => n1797);
   U73 : BUF_X1 port map( A => n1170, Z => n1785);
   U74 : BUF_X1 port map( A => n1155, Z => n1819);
   U75 : BUF_X1 port map( A => n1155, Z => n1818);
   U76 : BUF_X1 port map( A => n572, Z => n1906);
   U77 : BUF_X1 port map( A => n572, Z => n1905);
   U78 : BUF_X1 port map( A => n582, Z => n1882);
   U79 : BUF_X1 port map( A => n587, Z => n1870);
   U80 : BUF_X1 port map( A => n582, Z => n1881);
   U81 : BUF_X1 port map( A => n587, Z => n1869);
   U82 : BUF_X1 port map( A => n1138, Z => n1861);
   U83 : BUF_X1 port map( A => n1143, Z => n1849);
   U84 : BUF_X1 port map( A => n1148, Z => n1837);
   U85 : BUF_X1 port map( A => n1153, Z => n1825);
   U86 : BUF_X1 port map( A => n1163, Z => n1804);
   U87 : BUF_X1 port map( A => n1138, Z => n1860);
   U88 : BUF_X1 port map( A => n1143, Z => n1848);
   U89 : BUF_X1 port map( A => n1148, Z => n1836);
   U90 : BUF_X1 port map( A => n1153, Z => n1824);
   U91 : BUF_X1 port map( A => n1163, Z => n1803);
   U92 : BUF_X1 port map( A => n1166, Z => n1795);
   U93 : BUF_X1 port map( A => n1171, Z => n1783);
   U94 : BUF_X1 port map( A => n1166, Z => n1794);
   U95 : BUF_X1 port map( A => n1171, Z => n1782);
   U96 : BUF_X1 port map( A => n579, Z => n1889);
   U97 : BUF_X1 port map( A => n584, Z => n1877);
   U98 : BUF_X1 port map( A => n578, Z => n1891);
   U99 : BUF_X1 port map( A => n583, Z => n1879);
   U100 : BUF_X1 port map( A => n578, Z => n1890);
   U101 : BUF_X1 port map( A => n583, Z => n1878);
   U102 : BUF_X1 port map( A => n581, Z => n1885);
   U103 : BUF_X1 port map( A => n571, Z => n1909);
   U104 : BUF_X1 port map( A => n581, Z => n1884);
   U105 : BUF_X1 port map( A => n571, Z => n1908);
   U106 : BUF_X1 port map( A => n586, Z => n1873);
   U107 : BUF_X1 port map( A => n586, Z => n1872);
   U108 : BUF_X1 port map( A => n1160, Z => n1810);
   U109 : BUF_X1 port map( A => n1160, Z => n1809);
   U110 : BUF_X1 port map( A => n1135, Z => n1867);
   U111 : BUF_X1 port map( A => n1140, Z => n1855);
   U112 : BUF_X1 port map( A => n1145, Z => n1843);
   U113 : BUF_X1 port map( A => n1150, Z => n1831);
   U114 : BUF_X1 port map( A => n1135, Z => n1866);
   U115 : BUF_X1 port map( A => n1140, Z => n1854);
   U116 : BUF_X1 port map( A => n1145, Z => n1842);
   U117 : BUF_X1 port map( A => n1150, Z => n1830);
   U118 : BUF_X1 port map( A => n548, Z => n1961);
   U119 : BUF_X1 port map( A => n553, Z => n1949);
   U120 : BUF_X1 port map( A => n551, Z => n1955);
   U121 : BUF_X1 port map( A => n556, Z => n1943);
   U122 : BUF_X1 port map( A => n561, Z => n1931);
   U123 : BUF_X1 port map( A => n566, Z => n1919);
   U124 : BUF_X1 port map( A => n576, Z => n1898);
   U125 : BUF_X1 port map( A => n558, Z => n1937);
   U126 : BUF_X1 port map( A => n563, Z => n1925);
   U127 : BUF_X1 port map( A => n573, Z => n1904);
   U128 : BUF_X1 port map( A => n568, Z => n1913);
   U129 : BUF_X1 port map( A => n552, Z => n1952);
   U130 : BUF_X1 port map( A => n557, Z => n1940);
   U131 : BUF_X1 port map( A => n562, Z => n1928);
   U132 : BUF_X1 port map( A => n567, Z => n1916);
   U133 : BUF_X1 port map( A => n577, Z => n1895);
   U134 : BUF_X1 port map( A => n1158, Z => n1817);
   U135 : BUF_X1 port map( A => n1168, Z => n1793);
   U136 : BUF_X1 port map( A => n1173, Z => n1781);
   U137 : BUF_X1 port map( A => n1169, Z => n1790);
   U138 : BUF_X1 port map( A => n1174, Z => n1778);
   U139 : BUF_X1 port map( A => n1159, Z => n1814);
   U140 : BUF_X1 port map( A => n549, Z => n1957);
   U141 : BUF_X1 port map( A => n549, Z => n1956);
   U142 : BUF_X1 port map( A => n554, Z => n1945);
   U143 : BUF_X1 port map( A => n564, Z => n1921);
   U144 : BUF_X1 port map( A => n554, Z => n1944);
   U145 : BUF_X1 port map( A => n564, Z => n1920);
   U146 : BUF_X1 port map( A => n559, Z => n1933);
   U147 : BUF_X1 port map( A => n574, Z => n1900);
   U148 : BUF_X1 port map( A => n559, Z => n1932);
   U149 : BUF_X1 port map( A => n574, Z => n1899);
   U150 : BUF_X1 port map( A => n1139, Z => n1857);
   U151 : BUF_X1 port map( A => n1144, Z => n1845);
   U152 : BUF_X1 port map( A => n1149, Z => n1833);
   U153 : BUF_X1 port map( A => n1154, Z => n1821);
   U154 : BUF_X1 port map( A => n1164, Z => n1800);
   U155 : BUF_X1 port map( A => n1139, Z => n1858);
   U156 : BUF_X1 port map( A => n1144, Z => n1846);
   U157 : BUF_X1 port map( A => n1149, Z => n1834);
   U158 : BUF_X1 port map( A => n1154, Z => n1822);
   U159 : BUF_X1 port map( A => n1164, Z => n1801);
   U160 : BUF_X1 port map( A => n1161, Z => n1808);
   U161 : BUF_X1 port map( A => n1136, Z => n1865);
   U162 : BUF_X1 port map( A => n1141, Z => n1853);
   U163 : BUF_X1 port map( A => n1151, Z => n1829);
   U164 : BUF_X1 port map( A => n1146, Z => n1841);
   U165 : BUF_X1 port map( A => n1165, Z => n1799);
   U166 : BUF_X1 port map( A => n1170, Z => n1787);
   U167 : BUF_X1 port map( A => n1155, Z => n1820);
   U168 : BUF_X1 port map( A => n572, Z => n1907);
   U169 : BUF_X1 port map( A => n582, Z => n1883);
   U170 : BUF_X1 port map( A => n587, Z => n1871);
   U171 : BUF_X1 port map( A => n1138, Z => n1862);
   U172 : BUF_X1 port map( A => n1143, Z => n1850);
   U173 : BUF_X1 port map( A => n1148, Z => n1838);
   U174 : BUF_X1 port map( A => n1153, Z => n1826);
   U175 : BUF_X1 port map( A => n1163, Z => n1805);
   U176 : BUF_X1 port map( A => n1166, Z => n1796);
   U177 : BUF_X1 port map( A => n1171, Z => n1784);
   U178 : BUF_X1 port map( A => n578, Z => n1892);
   U179 : BUF_X1 port map( A => n583, Z => n1880);
   U180 : BUF_X1 port map( A => n581, Z => n1886);
   U181 : BUF_X1 port map( A => n571, Z => n1910);
   U182 : BUF_X1 port map( A => n586, Z => n1874);
   U183 : BUF_X1 port map( A => n1160, Z => n1811);
   U184 : BUF_X1 port map( A => n1135, Z => n1868);
   U185 : BUF_X1 port map( A => n1140, Z => n1856);
   U186 : BUF_X1 port map( A => n1145, Z => n1844);
   U187 : BUF_X1 port map( A => n1150, Z => n1832);
   U188 : BUF_X1 port map( A => n549, Z => n1958);
   U189 : BUF_X1 port map( A => n554, Z => n1946);
   U190 : BUF_X1 port map( A => n564, Z => n1922);
   U191 : BUF_X1 port map( A => n559, Z => n1934);
   U192 : BUF_X1 port map( A => n574, Z => n1901);
   U193 : BUF_X1 port map( A => n1139, Z => n1859);
   U194 : BUF_X1 port map( A => n1144, Z => n1847);
   U195 : BUF_X1 port map( A => n1149, Z => n1835);
   U196 : BUF_X1 port map( A => n1154, Z => n1823);
   U197 : BUF_X1 port map( A => n1164, Z => n1802);
   U198 : BUF_X1 port map( A => N307, Z => n2155);
   U199 : BUF_X1 port map( A => N307, Z => n2154);
   U200 : BUF_X1 port map( A => N340, Z => n2056);
   U201 : BUF_X1 port map( A => N340, Z => n2055);
   U202 : BUF_X1 port map( A => N341, Z => n2053);
   U203 : BUF_X1 port map( A => N341, Z => n2052);
   U204 : BUF_X1 port map( A => N342, Z => n2050);
   U205 : BUF_X1 port map( A => N342, Z => n2049);
   U206 : BUF_X1 port map( A => N343, Z => n2047);
   U207 : BUF_X1 port map( A => N343, Z => n2046);
   U208 : BUF_X1 port map( A => N344, Z => n2044);
   U209 : BUF_X1 port map( A => N344, Z => n2043);
   U210 : BUF_X1 port map( A => N345, Z => n2041);
   U211 : BUF_X1 port map( A => N345, Z => n2040);
   U212 : BUF_X1 port map( A => N346, Z => n2038);
   U213 : BUF_X1 port map( A => N346, Z => n2037);
   U214 : BUF_X1 port map( A => N347, Z => n2035);
   U215 : BUF_X1 port map( A => N347, Z => n2034);
   U216 : BUF_X1 port map( A => N348, Z => n2032);
   U217 : BUF_X1 port map( A => N348, Z => n2031);
   U218 : BUF_X1 port map( A => N349, Z => n2029);
   U219 : BUF_X1 port map( A => N349, Z => n2028);
   U220 : BUF_X1 port map( A => N350, Z => n2026);
   U221 : BUF_X1 port map( A => N350, Z => n2025);
   U222 : BUF_X1 port map( A => N351, Z => n2023);
   U223 : BUF_X1 port map( A => N351, Z => n2022);
   U224 : BUF_X1 port map( A => N352, Z => n2020);
   U225 : BUF_X1 port map( A => N352, Z => n2019);
   U226 : BUF_X1 port map( A => N353, Z => n2017);
   U227 : BUF_X1 port map( A => N353, Z => n2016);
   U228 : BUF_X1 port map( A => N354, Z => n2014);
   U229 : BUF_X1 port map( A => N354, Z => n2013);
   U230 : BUF_X1 port map( A => N355, Z => n2011);
   U231 : BUF_X1 port map( A => N355, Z => n2010);
   U232 : BUF_X1 port map( A => N356, Z => n2008);
   U233 : BUF_X1 port map( A => N356, Z => n2007);
   U234 : BUF_X1 port map( A => N357, Z => n2005);
   U235 : BUF_X1 port map( A => N357, Z => n2004);
   U236 : BUF_X1 port map( A => N358, Z => n2002);
   U237 : BUF_X1 port map( A => N358, Z => n2001);
   U238 : BUF_X1 port map( A => N359, Z => n1998);
   U239 : BUF_X1 port map( A => N359, Z => n1999);
   U240 : BUF_X1 port map( A => N360, Z => n1995);
   U241 : BUF_X1 port map( A => N360, Z => n1996);
   U242 : BUF_X1 port map( A => N361, Z => n1992);
   U243 : BUF_X1 port map( A => N361, Z => n1993);
   U244 : BUF_X1 port map( A => N362, Z => n1989);
   U245 : BUF_X1 port map( A => N362, Z => n1990);
   U246 : BUF_X1 port map( A => N363, Z => n1986);
   U247 : BUF_X1 port map( A => N363, Z => n1987);
   U248 : BUF_X1 port map( A => N364, Z => n1983);
   U249 : BUF_X1 port map( A => N364, Z => n1984);
   U250 : BUF_X1 port map( A => N365, Z => n1980);
   U251 : BUF_X1 port map( A => N365, Z => n1981);
   U252 : BUF_X1 port map( A => N366, Z => n1977);
   U253 : BUF_X1 port map( A => N366, Z => n1978);
   U254 : BUF_X1 port map( A => N367, Z => n1974);
   U255 : BUF_X1 port map( A => N367, Z => n1975);
   U256 : BUF_X1 port map( A => N368, Z => n1971);
   U257 : BUF_X1 port map( A => N368, Z => n1972);
   U258 : BUF_X1 port map( A => N369, Z => n1968);
   U259 : BUF_X1 port map( A => N369, Z => n1969);
   U260 : BUF_X1 port map( A => N308, Z => n2151);
   U261 : BUF_X1 port map( A => N316, Z => n2127);
   U262 : BUF_X1 port map( A => N317, Z => n2124);
   U263 : BUF_X1 port map( A => N318, Z => n2121);
   U264 : BUF_X1 port map( A => N319, Z => n2118);
   U265 : BUF_X1 port map( A => N320, Z => n2115);
   U266 : BUF_X1 port map( A => N321, Z => n2112);
   U267 : BUF_X1 port map( A => N322, Z => n2109);
   U268 : BUF_X1 port map( A => N323, Z => n2106);
   U269 : BUF_X1 port map( A => N324, Z => n2103);
   U270 : BUF_X1 port map( A => N325, Z => n2100);
   U271 : BUF_X1 port map( A => N326, Z => n2097);
   U272 : BUF_X1 port map( A => N327, Z => n2094);
   U273 : BUF_X1 port map( A => N328, Z => n2091);
   U274 : BUF_X1 port map( A => N329, Z => n2088);
   U275 : BUF_X1 port map( A => N330, Z => n2085);
   U276 : BUF_X1 port map( A => N331, Z => n2082);
   U277 : BUF_X1 port map( A => N332, Z => n2079);
   U278 : BUF_X1 port map( A => N333, Z => n2076);
   U279 : BUF_X1 port map( A => N334, Z => n2073);
   U280 : BUF_X1 port map( A => N335, Z => n2070);
   U281 : BUF_X1 port map( A => N336, Z => n2067);
   U282 : BUF_X1 port map( A => N337, Z => n2064);
   U283 : BUF_X1 port map( A => N338, Z => n2061);
   U284 : BUF_X1 port map( A => N339, Z => n2058);
   U285 : BUF_X1 port map( A => N308, Z => n2152);
   U286 : BUF_X1 port map( A => N316, Z => n2128);
   U287 : BUF_X1 port map( A => N317, Z => n2125);
   U288 : BUF_X1 port map( A => N318, Z => n2122);
   U289 : BUF_X1 port map( A => N319, Z => n2119);
   U290 : BUF_X1 port map( A => N320, Z => n2116);
   U291 : BUF_X1 port map( A => N321, Z => n2113);
   U292 : BUF_X1 port map( A => N322, Z => n2110);
   U293 : BUF_X1 port map( A => N323, Z => n2107);
   U294 : BUF_X1 port map( A => N324, Z => n2104);
   U295 : BUF_X1 port map( A => N325, Z => n2101);
   U296 : BUF_X1 port map( A => N326, Z => n2098);
   U297 : BUF_X1 port map( A => N327, Z => n2095);
   U298 : BUF_X1 port map( A => N328, Z => n2092);
   U299 : BUF_X1 port map( A => N329, Z => n2089);
   U300 : BUF_X1 port map( A => N330, Z => n2086);
   U301 : BUF_X1 port map( A => N331, Z => n2083);
   U302 : BUF_X1 port map( A => N332, Z => n2080);
   U303 : BUF_X1 port map( A => N333, Z => n2077);
   U304 : BUF_X1 port map( A => N334, Z => n2074);
   U305 : BUF_X1 port map( A => N335, Z => n2071);
   U306 : BUF_X1 port map( A => N336, Z => n2068);
   U307 : BUF_X1 port map( A => N337, Z => n2065);
   U308 : BUF_X1 port map( A => N338, Z => n2062);
   U309 : BUF_X1 port map( A => N339, Z => n2059);
   U310 : BUF_X1 port map( A => N309, Z => n2148);
   U311 : BUF_X1 port map( A => N310, Z => n2145);
   U312 : BUF_X1 port map( A => N311, Z => n2142);
   U313 : BUF_X1 port map( A => N312, Z => n2139);
   U314 : BUF_X1 port map( A => N313, Z => n2136);
   U315 : BUF_X1 port map( A => N314, Z => n2133);
   U316 : BUF_X1 port map( A => N315, Z => n2130);
   U317 : BUF_X1 port map( A => N309, Z => n2149);
   U318 : BUF_X1 port map( A => N310, Z => n2146);
   U319 : BUF_X1 port map( A => N311, Z => n2143);
   U320 : BUF_X1 port map( A => N312, Z => n2140);
   U321 : BUF_X1 port map( A => N313, Z => n2137);
   U322 : BUF_X1 port map( A => N314, Z => n2134);
   U323 : BUF_X1 port map( A => N315, Z => n2131);
   U324 : BUF_X1 port map( A => N307, Z => n2156);
   U325 : BUF_X1 port map( A => N340, Z => n2057);
   U326 : BUF_X1 port map( A => N341, Z => n2054);
   U327 : BUF_X1 port map( A => N342, Z => n2051);
   U328 : BUF_X1 port map( A => N343, Z => n2048);
   U329 : BUF_X1 port map( A => N344, Z => n2045);
   U330 : BUF_X1 port map( A => N345, Z => n2042);
   U331 : BUF_X1 port map( A => N346, Z => n2039);
   U332 : BUF_X1 port map( A => N347, Z => n2036);
   U333 : BUF_X1 port map( A => N348, Z => n2033);
   U334 : BUF_X1 port map( A => N349, Z => n2030);
   U335 : BUF_X1 port map( A => N350, Z => n2027);
   U336 : BUF_X1 port map( A => N351, Z => n2024);
   U337 : BUF_X1 port map( A => N352, Z => n2021);
   U338 : BUF_X1 port map( A => N353, Z => n2018);
   U339 : BUF_X1 port map( A => N354, Z => n2015);
   U340 : BUF_X1 port map( A => N355, Z => n2012);
   U341 : BUF_X1 port map( A => N356, Z => n2009);
   U342 : BUF_X1 port map( A => N357, Z => n2006);
   U343 : BUF_X1 port map( A => N358, Z => n2003);
   U344 : BUF_X1 port map( A => N359, Z => n2000);
   U345 : BUF_X1 port map( A => N360, Z => n1997);
   U346 : BUF_X1 port map( A => N361, Z => n1994);
   U347 : BUF_X1 port map( A => N362, Z => n1991);
   U348 : BUF_X1 port map( A => N363, Z => n1988);
   U349 : BUF_X1 port map( A => N364, Z => n1985);
   U350 : BUF_X1 port map( A => N365, Z => n1982);
   U351 : BUF_X1 port map( A => N366, Z => n1979);
   U352 : BUF_X1 port map( A => N367, Z => n1976);
   U353 : BUF_X1 port map( A => N368, Z => n1973);
   U354 : BUF_X1 port map( A => N369, Z => n1970);
   U355 : BUF_X1 port map( A => N308, Z => n2153);
   U356 : BUF_X1 port map( A => N316, Z => n2129);
   U357 : BUF_X1 port map( A => N317, Z => n2126);
   U358 : BUF_X1 port map( A => N318, Z => n2123);
   U359 : BUF_X1 port map( A => N319, Z => n2120);
   U360 : BUF_X1 port map( A => N320, Z => n2117);
   U361 : BUF_X1 port map( A => N321, Z => n2114);
   U362 : BUF_X1 port map( A => N322, Z => n2111);
   U363 : BUF_X1 port map( A => N323, Z => n2108);
   U364 : BUF_X1 port map( A => N324, Z => n2105);
   U365 : BUF_X1 port map( A => N325, Z => n2102);
   U366 : BUF_X1 port map( A => N326, Z => n2099);
   U367 : BUF_X1 port map( A => N327, Z => n2096);
   U368 : BUF_X1 port map( A => N328, Z => n2093);
   U369 : BUF_X1 port map( A => N329, Z => n2090);
   U370 : BUF_X1 port map( A => N330, Z => n2087);
   U371 : BUF_X1 port map( A => N331, Z => n2084);
   U372 : BUF_X1 port map( A => N332, Z => n2081);
   U373 : BUF_X1 port map( A => N333, Z => n2078);
   U374 : BUF_X1 port map( A => N334, Z => n2075);
   U375 : BUF_X1 port map( A => N335, Z => n2072);
   U376 : BUF_X1 port map( A => N336, Z => n2069);
   U377 : BUF_X1 port map( A => N337, Z => n2066);
   U378 : BUF_X1 port map( A => N338, Z => n2063);
   U379 : BUF_X1 port map( A => N339, Z => n2060);
   U380 : BUF_X1 port map( A => N309, Z => n2150);
   U381 : BUF_X1 port map( A => N310, Z => n2147);
   U382 : BUF_X1 port map( A => N311, Z => n2144);
   U383 : BUF_X1 port map( A => N312, Z => n2141);
   U384 : BUF_X1 port map( A => N313, Z => n2138);
   U385 : BUF_X1 port map( A => N314, Z => n2135);
   U386 : BUF_X1 port map( A => N315, Z => n2132);
   U387 : NOR2_X1 port map( A1 => n2683, A2 => n2682, ZN => n1699);
   U388 : NOR2_X1 port map( A1 => n2687, A2 => n2686, ZN => n1112);
   U389 : NOR4_X1 port map( A1 => n1298, A2 => n1299, A3 => n1300, A4 => n1301,
                           ZN => n1297);
   U390 : OAI221_X1 port map( B1 => n2672, B2 => n1831, C1 => n2640, C2 => 
                           n1828, A => n1305, ZN => n1298);
   U391 : OAI221_X1 port map( B1 => n2608, B2 => n1843, C1 => n2576, C2 => 
                           n1840, A => n1304, ZN => n1299);
   U392 : OAI221_X1 port map( B1 => n2544, B2 => n1855, C1 => n2512, C2 => 
                           n1852, A => n1303, ZN => n1300);
   U393 : NOR4_X1 port map( A1 => n1315, A2 => n1316, A3 => n1317, A4 => n1318,
                           ZN => n1314);
   U394 : OAI221_X1 port map( B1 => n2671, B2 => n1831, C1 => n2639, C2 => 
                           n1828, A => n1322, ZN => n1315);
   U395 : OAI221_X1 port map( B1 => n2607, B2 => n1843, C1 => n2575, C2 => 
                           n1840, A => n1321, ZN => n1316);
   U396 : OAI221_X1 port map( B1 => n2543, B2 => n1855, C1 => n2511, C2 => 
                           n1852, A => n1320, ZN => n1317);
   U397 : NOR4_X1 port map( A1 => n1332, A2 => n1333, A3 => n1334, A4 => n1335,
                           ZN => n1331);
   U398 : OAI221_X1 port map( B1 => n2670, B2 => n1831, C1 => n2638, C2 => 
                           n1828, A => n1339, ZN => n1332);
   U399 : OAI221_X1 port map( B1 => n2606, B2 => n1843, C1 => n2574, C2 => 
                           n1840, A => n1338, ZN => n1333);
   U400 : OAI221_X1 port map( B1 => n2542, B2 => n1855, C1 => n2510, C2 => 
                           n1852, A => n1337, ZN => n1334);
   U401 : NOR4_X1 port map( A1 => n1349, A2 => n1350, A3 => n1351, A4 => n1352,
                           ZN => n1348);
   U402 : OAI221_X1 port map( B1 => n2669, B2 => n1831, C1 => n2637, C2 => 
                           n1828, A => n1356, ZN => n1349);
   U403 : OAI221_X1 port map( B1 => n2605, B2 => n1843, C1 => n2573, C2 => 
                           n1840, A => n1355, ZN => n1350);
   U404 : OAI221_X1 port map( B1 => n2541, B2 => n1855, C1 => n2509, C2 => 
                           n1852, A => n1354, ZN => n1351);
   U405 : NOR4_X1 port map( A1 => n1366, A2 => n1367, A3 => n1368, A4 => n1369,
                           ZN => n1365);
   U406 : OAI221_X1 port map( B1 => n2668, B2 => n1831, C1 => n2636, C2 => 
                           n1828, A => n1373, ZN => n1366);
   U407 : OAI221_X1 port map( B1 => n2604, B2 => n1843, C1 => n2572, C2 => 
                           n1840, A => n1372, ZN => n1367);
   U408 : OAI221_X1 port map( B1 => n2540, B2 => n1855, C1 => n2508, C2 => 
                           n1852, A => n1371, ZN => n1368);
   U409 : NOR4_X1 port map( A1 => n1383, A2 => n1384, A3 => n1385, A4 => n1386,
                           ZN => n1382);
   U410 : OAI221_X1 port map( B1 => n2667, B2 => n1831, C1 => n2635, C2 => 
                           n1828, A => n1390, ZN => n1383);
   U411 : OAI221_X1 port map( B1 => n2603, B2 => n1843, C1 => n2571, C2 => 
                           n1840, A => n1389, ZN => n1384);
   U412 : OAI221_X1 port map( B1 => n2539, B2 => n1855, C1 => n2507, C2 => 
                           n1852, A => n1388, ZN => n1385);
   U413 : NOR4_X1 port map( A1 => n1400, A2 => n1401, A3 => n1402, A4 => n1403,
                           ZN => n1399);
   U414 : OAI221_X1 port map( B1 => n2666, B2 => n1831, C1 => n2634, C2 => 
                           n1828, A => n1407, ZN => n1400);
   U415 : OAI221_X1 port map( B1 => n2602, B2 => n1843, C1 => n2570, C2 => 
                           n1840, A => n1406, ZN => n1401);
   U416 : OAI221_X1 port map( B1 => n2538, B2 => n1855, C1 => n2506, C2 => 
                           n1852, A => n1405, ZN => n1402);
   U417 : NOR4_X1 port map( A1 => n1417, A2 => n1418, A3 => n1419, A4 => n1420,
                           ZN => n1416);
   U418 : OAI221_X1 port map( B1 => n2665, B2 => n1831, C1 => n2633, C2 => 
                           n1828, A => n1424, ZN => n1417);
   U419 : OAI221_X1 port map( B1 => n2601, B2 => n1843, C1 => n2569, C2 => 
                           n1840, A => n1423, ZN => n1418);
   U420 : OAI221_X1 port map( B1 => n2537, B2 => n1855, C1 => n2505, C2 => 
                           n1852, A => n1422, ZN => n1419);
   U421 : NOR4_X1 port map( A1 => n1434, A2 => n1435, A3 => n1436, A4 => n1437,
                           ZN => n1433);
   U422 : OAI221_X1 port map( B1 => n2664, B2 => n1831, C1 => n2632, C2 => 
                           n1828, A => n1441, ZN => n1434);
   U423 : OAI221_X1 port map( B1 => n2600, B2 => n1843, C1 => n2568, C2 => 
                           n1840, A => n1440, ZN => n1435);
   U424 : OAI221_X1 port map( B1 => n2536, B2 => n1855, C1 => n2504, C2 => 
                           n1852, A => n1439, ZN => n1436);
   U425 : NOR4_X1 port map( A1 => n1451, A2 => n1452, A3 => n1453, A4 => n1454,
                           ZN => n1450);
   U426 : OAI221_X1 port map( B1 => n2663, B2 => n1831, C1 => n2631, C2 => 
                           n1828, A => n1458, ZN => n1451);
   U427 : OAI221_X1 port map( B1 => n2599, B2 => n1843, C1 => n2567, C2 => 
                           n1840, A => n1457, ZN => n1452);
   U428 : OAI221_X1 port map( B1 => n2535, B2 => n1855, C1 => n2503, C2 => 
                           n1852, A => n1456, ZN => n1453);
   U429 : NOR4_X1 port map( A1 => n1468, A2 => n1469, A3 => n1470, A4 => n1471,
                           ZN => n1467);
   U430 : OAI221_X1 port map( B1 => n2662, B2 => n1831, C1 => n2630, C2 => 
                           n1828, A => n1475, ZN => n1468);
   U431 : OAI221_X1 port map( B1 => n2598, B2 => n1843, C1 => n2566, C2 => 
                           n1840, A => n1474, ZN => n1469);
   U432 : OAI221_X1 port map( B1 => n2534, B2 => n1855, C1 => n2502, C2 => 
                           n1852, A => n1473, ZN => n1470);
   U433 : NOR4_X1 port map( A1 => n1485, A2 => n1486, A3 => n1487, A4 => n1488,
                           ZN => n1484);
   U434 : OAI221_X1 port map( B1 => n2661, B2 => n1831, C1 => n2629, C2 => 
                           n1828, A => n1492, ZN => n1485);
   U435 : OAI221_X1 port map( B1 => n2597, B2 => n1843, C1 => n2565, C2 => 
                           n1840, A => n1491, ZN => n1486);
   U436 : OAI221_X1 port map( B1 => n2533, B2 => n1855, C1 => n2501, C2 => 
                           n1852, A => n1490, ZN => n1487);
   U437 : NOR4_X1 port map( A1 => n1502, A2 => n1503, A3 => n1504, A4 => n1505,
                           ZN => n1501);
   U438 : OAI221_X1 port map( B1 => n2660, B2 => n1830, C1 => n2628, C2 => 
                           n1827, A => n1509, ZN => n1502);
   U439 : OAI221_X1 port map( B1 => n2596, B2 => n1842, C1 => n2564, C2 => 
                           n1839, A => n1508, ZN => n1503);
   U440 : OAI221_X1 port map( B1 => n2532, B2 => n1854, C1 => n2500, C2 => 
                           n1851, A => n1507, ZN => n1504);
   U441 : NOR4_X1 port map( A1 => n1519, A2 => n1520, A3 => n1521, A4 => n1522,
                           ZN => n1518);
   U442 : OAI221_X1 port map( B1 => n2659, B2 => n1830, C1 => n2627, C2 => 
                           n1827, A => n1526, ZN => n1519);
   U443 : OAI221_X1 port map( B1 => n2595, B2 => n1842, C1 => n2563, C2 => 
                           n1839, A => n1525, ZN => n1520);
   U444 : OAI221_X1 port map( B1 => n2531, B2 => n1854, C1 => n2499, C2 => 
                           n1851, A => n1524, ZN => n1521);
   U445 : NOR4_X1 port map( A1 => n1536, A2 => n1537, A3 => n1538, A4 => n1539,
                           ZN => n1535);
   U446 : OAI221_X1 port map( B1 => n2658, B2 => n1830, C1 => n2626, C2 => 
                           n1827, A => n1543, ZN => n1536);
   U447 : OAI221_X1 port map( B1 => n2594, B2 => n1842, C1 => n2562, C2 => 
                           n1839, A => n1542, ZN => n1537);
   U448 : OAI221_X1 port map( B1 => n2530, B2 => n1854, C1 => n2498, C2 => 
                           n1851, A => n1541, ZN => n1538);
   U449 : NOR4_X1 port map( A1 => n1553, A2 => n1554, A3 => n1555, A4 => n1556,
                           ZN => n1552);
   U450 : OAI221_X1 port map( B1 => n2657, B2 => n1830, C1 => n2625, C2 => 
                           n1827, A => n1560, ZN => n1553);
   U451 : OAI221_X1 port map( B1 => n2593, B2 => n1842, C1 => n2561, C2 => 
                           n1839, A => n1559, ZN => n1554);
   U452 : OAI221_X1 port map( B1 => n2529, B2 => n1854, C1 => n2497, C2 => 
                           n1851, A => n1558, ZN => n1555);
   U453 : NOR4_X1 port map( A1 => n1570, A2 => n1571, A3 => n1572, A4 => n1573,
                           ZN => n1569);
   U454 : OAI221_X1 port map( B1 => n2656, B2 => n1830, C1 => n2624, C2 => 
                           n1827, A => n1577, ZN => n1570);
   U455 : OAI221_X1 port map( B1 => n2592, B2 => n1842, C1 => n2560, C2 => 
                           n1839, A => n1576, ZN => n1571);
   U456 : OAI221_X1 port map( B1 => n2528, B2 => n1854, C1 => n2496, C2 => 
                           n1851, A => n1575, ZN => n1572);
   U457 : NOR4_X1 port map( A1 => n1587, A2 => n1588, A3 => n1589, A4 => n1590,
                           ZN => n1586);
   U458 : OAI221_X1 port map( B1 => n2655, B2 => n1830, C1 => n2623, C2 => 
                           n1827, A => n1594, ZN => n1587);
   U459 : OAI221_X1 port map( B1 => n2591, B2 => n1842, C1 => n2559, C2 => 
                           n1839, A => n1593, ZN => n1588);
   U460 : OAI221_X1 port map( B1 => n2527, B2 => n1854, C1 => n2495, C2 => 
                           n1851, A => n1592, ZN => n1589);
   U461 : NOR4_X1 port map( A1 => n1604, A2 => n1605, A3 => n1606, A4 => n1607,
                           ZN => n1603);
   U462 : OAI221_X1 port map( B1 => n2654, B2 => n1830, C1 => n2622, C2 => 
                           n1827, A => n1611, ZN => n1604);
   U463 : OAI221_X1 port map( B1 => n2590, B2 => n1842, C1 => n2558, C2 => 
                           n1839, A => n1610, ZN => n1605);
   U464 : OAI221_X1 port map( B1 => n2526, B2 => n1854, C1 => n2494, C2 => 
                           n1851, A => n1609, ZN => n1606);
   U465 : NOR4_X1 port map( A1 => n1621, A2 => n1622, A3 => n1623, A4 => n1624,
                           ZN => n1620);
   U466 : OAI221_X1 port map( B1 => n2653, B2 => n1830, C1 => n2621, C2 => 
                           n1827, A => n1628, ZN => n1621);
   U467 : OAI221_X1 port map( B1 => n2589, B2 => n1842, C1 => n2557, C2 => 
                           n1839, A => n1627, ZN => n1622);
   U468 : OAI221_X1 port map( B1 => n2525, B2 => n1854, C1 => n2493, C2 => 
                           n1851, A => n1626, ZN => n1623);
   U469 : NOR4_X1 port map( A1 => n1638, A2 => n1639, A3 => n1640, A4 => n1641,
                           ZN => n1637);
   U470 : OAI221_X1 port map( B1 => n2652, B2 => n1830, C1 => n2620, C2 => 
                           n1827, A => n1645, ZN => n1638);
   U471 : OAI221_X1 port map( B1 => n2588, B2 => n1842, C1 => n2556, C2 => 
                           n1839, A => n1644, ZN => n1639);
   U472 : OAI221_X1 port map( B1 => n2524, B2 => n1854, C1 => n2492, C2 => 
                           n1851, A => n1643, ZN => n1640);
   U473 : NOR4_X1 port map( A1 => n1655, A2 => n1656, A3 => n1657, A4 => n1658,
                           ZN => n1654);
   U474 : OAI221_X1 port map( B1 => n2651, B2 => n1830, C1 => n2619, C2 => 
                           n1827, A => n1662, ZN => n1655);
   U475 : OAI221_X1 port map( B1 => n2587, B2 => n1842, C1 => n2555, C2 => 
                           n1839, A => n1661, ZN => n1656);
   U476 : OAI221_X1 port map( B1 => n2523, B2 => n1854, C1 => n2491, C2 => 
                           n1851, A => n1660, ZN => n1657);
   U477 : NOR4_X1 port map( A1 => n1672, A2 => n1673, A3 => n1674, A4 => n1675,
                           ZN => n1671);
   U478 : OAI221_X1 port map( B1 => n2650, B2 => n1830, C1 => n2618, C2 => 
                           n1827, A => n1679, ZN => n1672);
   U479 : OAI221_X1 port map( B1 => n2586, B2 => n1842, C1 => n2554, C2 => 
                           n1839, A => n1678, ZN => n1673);
   U480 : OAI221_X1 port map( B1 => n2522, B2 => n1854, C1 => n2490, C2 => 
                           n1851, A => n1677, ZN => n1674);
   U481 : NOR4_X1 port map( A1 => n1689, A2 => n1690, A3 => n1691, A4 => n1692,
                           ZN => n1688);
   U482 : OAI221_X1 port map( B1 => n2649, B2 => n1830, C1 => n2617, C2 => 
                           n1827, A => n1704, ZN => n1689);
   U483 : OAI221_X1 port map( B1 => n2585, B2 => n1842, C1 => n2553, C2 => 
                           n1839, A => n1701, ZN => n1690);
   U484 : OAI221_X1 port map( B1 => n2521, B2 => n1854, C1 => n2489, C2 => 
                           n1851, A => n1698, ZN => n1691);
   U485 : NOR4_X1 port map( A1 => n1131, A2 => n1132, A3 => n1133, A4 => n1134,
                           ZN => n1130);
   U486 : OAI221_X1 port map( B1 => n2680, B2 => n1832, C1 => n2648, C2 => 
                           n1829, A => n1152, ZN => n1131);
   U487 : OAI221_X1 port map( B1 => n2616, B2 => n1844, C1 => n2584, C2 => 
                           n1841, A => n1147, ZN => n1132);
   U488 : OAI221_X1 port map( B1 => n2552, B2 => n1856, C1 => n2520, C2 => 
                           n1853, A => n1142, ZN => n1133);
   U489 : NOR4_X1 port map( A1 => n1179, A2 => n1180, A3 => n1181, A4 => n1182,
                           ZN => n1178);
   U490 : OAI221_X1 port map( B1 => n2679, B2 => n1832, C1 => n2647, C2 => 
                           n1829, A => n1186, ZN => n1179);
   U491 : OAI221_X1 port map( B1 => n2615, B2 => n1844, C1 => n2583, C2 => 
                           n1841, A => n1185, ZN => n1180);
   U492 : OAI221_X1 port map( B1 => n2551, B2 => n1856, C1 => n2519, C2 => 
                           n1853, A => n1184, ZN => n1181);
   U493 : NOR4_X1 port map( A1 => n1196, A2 => n1197, A3 => n1198, A4 => n1199,
                           ZN => n1195);
   U494 : OAI221_X1 port map( B1 => n2678, B2 => n1832, C1 => n2646, C2 => 
                           n1829, A => n1203, ZN => n1196);
   U495 : OAI221_X1 port map( B1 => n2614, B2 => n1844, C1 => n2582, C2 => 
                           n1841, A => n1202, ZN => n1197);
   U496 : OAI221_X1 port map( B1 => n2550, B2 => n1856, C1 => n2518, C2 => 
                           n1853, A => n1201, ZN => n1198);
   U497 : NOR4_X1 port map( A1 => n1213, A2 => n1214, A3 => n1215, A4 => n1216,
                           ZN => n1212);
   U498 : OAI221_X1 port map( B1 => n2677, B2 => n1832, C1 => n2645, C2 => 
                           n1829, A => n1220, ZN => n1213);
   U499 : OAI221_X1 port map( B1 => n2613, B2 => n1844, C1 => n2581, C2 => 
                           n1841, A => n1219, ZN => n1214);
   U500 : OAI221_X1 port map( B1 => n2549, B2 => n1856, C1 => n2517, C2 => 
                           n1853, A => n1218, ZN => n1215);
   U501 : NOR4_X1 port map( A1 => n1230, A2 => n1231, A3 => n1232, A4 => n1233,
                           ZN => n1229);
   U502 : OAI221_X1 port map( B1 => n2676, B2 => n1832, C1 => n2644, C2 => 
                           n1829, A => n1237, ZN => n1230);
   U503 : OAI221_X1 port map( B1 => n2612, B2 => n1844, C1 => n2580, C2 => 
                           n1841, A => n1236, ZN => n1231);
   U504 : OAI221_X1 port map( B1 => n2548, B2 => n1856, C1 => n2516, C2 => 
                           n1853, A => n1235, ZN => n1232);
   U505 : NOR4_X1 port map( A1 => n1247, A2 => n1248, A3 => n1249, A4 => n1250,
                           ZN => n1246);
   U506 : OAI221_X1 port map( B1 => n2675, B2 => n1832, C1 => n2643, C2 => 
                           n1829, A => n1254, ZN => n1247);
   U507 : OAI221_X1 port map( B1 => n2611, B2 => n1844, C1 => n2579, C2 => 
                           n1841, A => n1253, ZN => n1248);
   U508 : OAI221_X1 port map( B1 => n2547, B2 => n1856, C1 => n2515, C2 => 
                           n1853, A => n1252, ZN => n1249);
   U509 : NOR4_X1 port map( A1 => n1264, A2 => n1265, A3 => n1266, A4 => n1267,
                           ZN => n1263);
   U510 : OAI221_X1 port map( B1 => n2674, B2 => n1832, C1 => n2642, C2 => 
                           n1829, A => n1271, ZN => n1264);
   U511 : OAI221_X1 port map( B1 => n2610, B2 => n1844, C1 => n2578, C2 => 
                           n1841, A => n1270, ZN => n1265);
   U512 : OAI221_X1 port map( B1 => n2546, B2 => n1856, C1 => n2514, C2 => 
                           n1853, A => n1269, ZN => n1266);
   U513 : NOR4_X1 port map( A1 => n1281, A2 => n1282, A3 => n1283, A4 => n1284,
                           ZN => n1280);
   U514 : OAI221_X1 port map( B1 => n2673, B2 => n1832, C1 => n2641, C2 => 
                           n1829, A => n1288, ZN => n1281);
   U515 : OAI221_X1 port map( B1 => n2609, B2 => n1844, C1 => n2577, C2 => 
                           n1841, A => n1287, ZN => n1282);
   U516 : OAI221_X1 port map( B1 => n2545, B2 => n1856, C1 => n2513, C2 => 
                           n1853, A => n1286, ZN => n1283);
   U517 : NOR4_X1 port map( A1 => n544, A2 => n545, A3 => n546, A4 => n547, ZN 
                           => n543);
   U518 : OAI221_X1 port map( B1 => n1925, B2 => n2680, C1 => n1922, C2 => 
                           n2648, A => n565, ZN => n544);
   U519 : OAI221_X1 port map( B1 => n1937, B2 => n2616, C1 => n1934, C2 => 
                           n2584, A => n560, ZN => n545);
   U520 : OAI221_X1 port map( B1 => n1949, B2 => n2552, C1 => n1946, C2 => 
                           n2520, A => n555, ZN => n546);
   U521 : NOR4_X1 port map( A1 => n592, A2 => n593, A3 => n594, A4 => n595, ZN 
                           => n591);
   U522 : OAI221_X1 port map( B1 => n1925, B2 => n2679, C1 => n1922, C2 => 
                           n2647, A => n599, ZN => n592);
   U523 : OAI221_X1 port map( B1 => n1937, B2 => n2615, C1 => n1934, C2 => 
                           n2583, A => n598, ZN => n593);
   U524 : OAI221_X1 port map( B1 => n1949, B2 => n2551, C1 => n1946, C2 => 
                           n2519, A => n597, ZN => n594);
   U525 : NOR4_X1 port map( A1 => n609, A2 => n610, A3 => n611, A4 => n612, ZN 
                           => n608);
   U526 : OAI221_X1 port map( B1 => n1925, B2 => n2678, C1 => n1922, C2 => 
                           n2646, A => n616, ZN => n609);
   U527 : OAI221_X1 port map( B1 => n1937, B2 => n2614, C1 => n1934, C2 => 
                           n2582, A => n615, ZN => n610);
   U528 : OAI221_X1 port map( B1 => n1949, B2 => n2550, C1 => n1946, C2 => 
                           n2518, A => n614, ZN => n611);
   U529 : NOR4_X1 port map( A1 => n626, A2 => n627, A3 => n628, A4 => n629, ZN 
                           => n625);
   U530 : OAI221_X1 port map( B1 => n1925, B2 => n2677, C1 => n1922, C2 => 
                           n2645, A => n633, ZN => n626);
   U531 : OAI221_X1 port map( B1 => n1937, B2 => n2613, C1 => n1934, C2 => 
                           n2581, A => n632, ZN => n627);
   U532 : OAI221_X1 port map( B1 => n1949, B2 => n2549, C1 => n1946, C2 => 
                           n2517, A => n631, ZN => n628);
   U533 : NOR4_X1 port map( A1 => n643, A2 => n644, A3 => n645, A4 => n646, ZN 
                           => n642);
   U534 : OAI221_X1 port map( B1 => n1925, B2 => n2676, C1 => n1922, C2 => 
                           n2644, A => n650, ZN => n643);
   U535 : OAI221_X1 port map( B1 => n1937, B2 => n2612, C1 => n1934, C2 => 
                           n2580, A => n649, ZN => n644);
   U536 : OAI221_X1 port map( B1 => n1949, B2 => n2548, C1 => n1946, C2 => 
                           n2516, A => n648, ZN => n645);
   U537 : NOR4_X1 port map( A1 => n660, A2 => n661, A3 => n662, A4 => n663, ZN 
                           => n659);
   U538 : OAI221_X1 port map( B1 => n1925, B2 => n2675, C1 => n1922, C2 => 
                           n2643, A => n667, ZN => n660);
   U539 : OAI221_X1 port map( B1 => n1937, B2 => n2611, C1 => n1934, C2 => 
                           n2579, A => n666, ZN => n661);
   U540 : OAI221_X1 port map( B1 => n1949, B2 => n2547, C1 => n1946, C2 => 
                           n2515, A => n665, ZN => n662);
   U541 : NOR4_X1 port map( A1 => n677, A2 => n678, A3 => n679, A4 => n680, ZN 
                           => n676);
   U542 : OAI221_X1 port map( B1 => n1925, B2 => n2674, C1 => n1922, C2 => 
                           n2642, A => n684, ZN => n677);
   U543 : OAI221_X1 port map( B1 => n1937, B2 => n2610, C1 => n1934, C2 => 
                           n2578, A => n683, ZN => n678);
   U544 : OAI221_X1 port map( B1 => n1949, B2 => n2546, C1 => n1946, C2 => 
                           n2514, A => n682, ZN => n679);
   U545 : NOR4_X1 port map( A1 => n694, A2 => n695, A3 => n696, A4 => n697, ZN 
                           => n693);
   U546 : OAI221_X1 port map( B1 => n1925, B2 => n2673, C1 => n1922, C2 => 
                           n2641, A => n701, ZN => n694);
   U547 : OAI221_X1 port map( B1 => n1937, B2 => n2609, C1 => n1934, C2 => 
                           n2577, A => n700, ZN => n695);
   U548 : OAI221_X1 port map( B1 => n1949, B2 => n2545, C1 => n1946, C2 => 
                           n2513, A => n699, ZN => n696);
   U549 : NOR4_X1 port map( A1 => n711, A2 => n712, A3 => n713, A4 => n714, ZN 
                           => n710);
   U550 : OAI221_X1 port map( B1 => n1924, B2 => n2672, C1 => n1921, C2 => 
                           n2640, A => n718, ZN => n711);
   U551 : OAI221_X1 port map( B1 => n1936, B2 => n2608, C1 => n1933, C2 => 
                           n2576, A => n717, ZN => n712);
   U552 : OAI221_X1 port map( B1 => n1948, B2 => n2544, C1 => n1945, C2 => 
                           n2512, A => n716, ZN => n713);
   U553 : NOR4_X1 port map( A1 => n728, A2 => n729, A3 => n730, A4 => n731, ZN 
                           => n727);
   U554 : OAI221_X1 port map( B1 => n1924, B2 => n2671, C1 => n1921, C2 => 
                           n2639, A => n735, ZN => n728);
   U555 : OAI221_X1 port map( B1 => n1936, B2 => n2607, C1 => n1933, C2 => 
                           n2575, A => n734, ZN => n729);
   U556 : OAI221_X1 port map( B1 => n1948, B2 => n2543, C1 => n1945, C2 => 
                           n2511, A => n733, ZN => n730);
   U557 : NOR4_X1 port map( A1 => n745, A2 => n746, A3 => n747, A4 => n748, ZN 
                           => n744);
   U558 : OAI221_X1 port map( B1 => n1924, B2 => n2670, C1 => n1921, C2 => 
                           n2638, A => n752, ZN => n745);
   U559 : OAI221_X1 port map( B1 => n1936, B2 => n2606, C1 => n1933, C2 => 
                           n2574, A => n751, ZN => n746);
   U560 : OAI221_X1 port map( B1 => n1948, B2 => n2542, C1 => n1945, C2 => 
                           n2510, A => n750, ZN => n747);
   U561 : NOR4_X1 port map( A1 => n762, A2 => n763, A3 => n764, A4 => n765, ZN 
                           => n761);
   U562 : OAI221_X1 port map( B1 => n1924, B2 => n2669, C1 => n1921, C2 => 
                           n2637, A => n769, ZN => n762);
   U563 : OAI221_X1 port map( B1 => n1936, B2 => n2605, C1 => n1933, C2 => 
                           n2573, A => n768, ZN => n763);
   U564 : OAI221_X1 port map( B1 => n1948, B2 => n2541, C1 => n1945, C2 => 
                           n2509, A => n767, ZN => n764);
   U565 : NOR4_X1 port map( A1 => n779, A2 => n780, A3 => n781, A4 => n782, ZN 
                           => n778);
   U566 : OAI221_X1 port map( B1 => n1924, B2 => n2668, C1 => n1921, C2 => 
                           n2636, A => n786, ZN => n779);
   U567 : OAI221_X1 port map( B1 => n1936, B2 => n2604, C1 => n1933, C2 => 
                           n2572, A => n785, ZN => n780);
   U568 : OAI221_X1 port map( B1 => n1948, B2 => n2540, C1 => n1945, C2 => 
                           n2508, A => n784, ZN => n781);
   U569 : NOR4_X1 port map( A1 => n796, A2 => n797, A3 => n798, A4 => n799, ZN 
                           => n795);
   U570 : OAI221_X1 port map( B1 => n1924, B2 => n2667, C1 => n1921, C2 => 
                           n2635, A => n803, ZN => n796);
   U571 : OAI221_X1 port map( B1 => n1936, B2 => n2603, C1 => n1933, C2 => 
                           n2571, A => n802, ZN => n797);
   U572 : OAI221_X1 port map( B1 => n1948, B2 => n2539, C1 => n1945, C2 => 
                           n2507, A => n801, ZN => n798);
   U573 : NOR4_X1 port map( A1 => n813, A2 => n814, A3 => n815, A4 => n816, ZN 
                           => n812);
   U574 : OAI221_X1 port map( B1 => n1924, B2 => n2666, C1 => n1921, C2 => 
                           n2634, A => n820, ZN => n813);
   U575 : OAI221_X1 port map( B1 => n1936, B2 => n2602, C1 => n1933, C2 => 
                           n2570, A => n819, ZN => n814);
   U576 : OAI221_X1 port map( B1 => n1948, B2 => n2538, C1 => n1945, C2 => 
                           n2506, A => n818, ZN => n815);
   U577 : NOR4_X1 port map( A1 => n830, A2 => n831, A3 => n832, A4 => n833, ZN 
                           => n829);
   U578 : OAI221_X1 port map( B1 => n1924, B2 => n2665, C1 => n1921, C2 => 
                           n2633, A => n837, ZN => n830);
   U579 : OAI221_X1 port map( B1 => n1936, B2 => n2601, C1 => n1933, C2 => 
                           n2569, A => n836, ZN => n831);
   U580 : OAI221_X1 port map( B1 => n1948, B2 => n2537, C1 => n1945, C2 => 
                           n2505, A => n835, ZN => n832);
   U581 : NOR4_X1 port map( A1 => n847, A2 => n848, A3 => n849, A4 => n850, ZN 
                           => n846);
   U582 : OAI221_X1 port map( B1 => n1924, B2 => n2664, C1 => n1921, C2 => 
                           n2632, A => n854, ZN => n847);
   U583 : OAI221_X1 port map( B1 => n1936, B2 => n2600, C1 => n1933, C2 => 
                           n2568, A => n853, ZN => n848);
   U584 : OAI221_X1 port map( B1 => n1948, B2 => n2536, C1 => n1945, C2 => 
                           n2504, A => n852, ZN => n849);
   U585 : NOR4_X1 port map( A1 => n864, A2 => n865, A3 => n866, A4 => n867, ZN 
                           => n863);
   U586 : OAI221_X1 port map( B1 => n1924, B2 => n2663, C1 => n1921, C2 => 
                           n2631, A => n871, ZN => n864);
   U587 : OAI221_X1 port map( B1 => n1936, B2 => n2599, C1 => n1933, C2 => 
                           n2567, A => n870, ZN => n865);
   U588 : OAI221_X1 port map( B1 => n1948, B2 => n2535, C1 => n1945, C2 => 
                           n2503, A => n869, ZN => n866);
   U589 : NOR4_X1 port map( A1 => n881, A2 => n882, A3 => n883, A4 => n884, ZN 
                           => n880);
   U590 : OAI221_X1 port map( B1 => n1924, B2 => n2662, C1 => n1921, C2 => 
                           n2630, A => n888, ZN => n881);
   U591 : OAI221_X1 port map( B1 => n1936, B2 => n2598, C1 => n1933, C2 => 
                           n2566, A => n887, ZN => n882);
   U592 : OAI221_X1 port map( B1 => n1948, B2 => n2534, C1 => n1945, C2 => 
                           n2502, A => n886, ZN => n883);
   U593 : NOR4_X1 port map( A1 => n898, A2 => n899, A3 => n900, A4 => n901, ZN 
                           => n897);
   U594 : OAI221_X1 port map( B1 => n1924, B2 => n2661, C1 => n1921, C2 => 
                           n2629, A => n905, ZN => n898);
   U595 : OAI221_X1 port map( B1 => n1936, B2 => n2597, C1 => n1933, C2 => 
                           n2565, A => n904, ZN => n899);
   U596 : OAI221_X1 port map( B1 => n1948, B2 => n2533, C1 => n1945, C2 => 
                           n2501, A => n903, ZN => n900);
   U597 : NOR4_X1 port map( A1 => n915, A2 => n916, A3 => n917, A4 => n918, ZN 
                           => n914);
   U598 : OAI221_X1 port map( B1 => n1923, B2 => n2660, C1 => n1920, C2 => 
                           n2628, A => n922, ZN => n915);
   U599 : OAI221_X1 port map( B1 => n1935, B2 => n2596, C1 => n1932, C2 => 
                           n2564, A => n921, ZN => n916);
   U600 : OAI221_X1 port map( B1 => n1947, B2 => n2532, C1 => n1944, C2 => 
                           n2500, A => n920, ZN => n917);
   U601 : NOR4_X1 port map( A1 => n932, A2 => n933, A3 => n934, A4 => n935, ZN 
                           => n931);
   U602 : OAI221_X1 port map( B1 => n1923, B2 => n2659, C1 => n1920, C2 => 
                           n2627, A => n939, ZN => n932);
   U603 : OAI221_X1 port map( B1 => n1935, B2 => n2595, C1 => n1932, C2 => 
                           n2563, A => n938, ZN => n933);
   U604 : OAI221_X1 port map( B1 => n1947, B2 => n2531, C1 => n1944, C2 => 
                           n2499, A => n937, ZN => n934);
   U605 : NOR4_X1 port map( A1 => n949, A2 => n950, A3 => n951, A4 => n952, ZN 
                           => n948);
   U606 : OAI221_X1 port map( B1 => n1923, B2 => n2658, C1 => n1920, C2 => 
                           n2626, A => n956, ZN => n949);
   U607 : OAI221_X1 port map( B1 => n1935, B2 => n2594, C1 => n1932, C2 => 
                           n2562, A => n955, ZN => n950);
   U608 : OAI221_X1 port map( B1 => n1947, B2 => n2530, C1 => n1944, C2 => 
                           n2498, A => n954, ZN => n951);
   U609 : NOR4_X1 port map( A1 => n966, A2 => n967, A3 => n968, A4 => n969, ZN 
                           => n965);
   U610 : OAI221_X1 port map( B1 => n1923, B2 => n2657, C1 => n1920, C2 => 
                           n2625, A => n973, ZN => n966);
   U611 : OAI221_X1 port map( B1 => n1935, B2 => n2593, C1 => n1932, C2 => 
                           n2561, A => n972, ZN => n967);
   U612 : OAI221_X1 port map( B1 => n1947, B2 => n2529, C1 => n1944, C2 => 
                           n2497, A => n971, ZN => n968);
   U613 : NOR4_X1 port map( A1 => n983, A2 => n984, A3 => n985, A4 => n986, ZN 
                           => n982);
   U614 : OAI221_X1 port map( B1 => n1923, B2 => n2656, C1 => n1920, C2 => 
                           n2624, A => n990, ZN => n983);
   U615 : OAI221_X1 port map( B1 => n1935, B2 => n2592, C1 => n1932, C2 => 
                           n2560, A => n989, ZN => n984);
   U616 : OAI221_X1 port map( B1 => n1947, B2 => n2528, C1 => n1944, C2 => 
                           n2496, A => n988, ZN => n985);
   U617 : NOR4_X1 port map( A1 => n1000, A2 => n1001, A3 => n1002, A4 => n1003,
                           ZN => n999);
   U618 : OAI221_X1 port map( B1 => n1923, B2 => n2655, C1 => n1920, C2 => 
                           n2623, A => n1007, ZN => n1000);
   U619 : OAI221_X1 port map( B1 => n1935, B2 => n2591, C1 => n1932, C2 => 
                           n2559, A => n1006, ZN => n1001);
   U620 : OAI221_X1 port map( B1 => n1947, B2 => n2527, C1 => n1944, C2 => 
                           n2495, A => n1005, ZN => n1002);
   U621 : NOR4_X1 port map( A1 => n1017, A2 => n1018, A3 => n1019, A4 => n1020,
                           ZN => n1016);
   U622 : OAI221_X1 port map( B1 => n1923, B2 => n2654, C1 => n1920, C2 => 
                           n2622, A => n1024, ZN => n1017);
   U623 : OAI221_X1 port map( B1 => n1935, B2 => n2590, C1 => n1932, C2 => 
                           n2558, A => n1023, ZN => n1018);
   U624 : OAI221_X1 port map( B1 => n1947, B2 => n2526, C1 => n1944, C2 => 
                           n2494, A => n1022, ZN => n1019);
   U625 : NOR4_X1 port map( A1 => n1034, A2 => n1035, A3 => n1036, A4 => n1037,
                           ZN => n1033);
   U626 : OAI221_X1 port map( B1 => n1923, B2 => n2653, C1 => n1920, C2 => 
                           n2621, A => n1041, ZN => n1034);
   U627 : OAI221_X1 port map( B1 => n1935, B2 => n2589, C1 => n1932, C2 => 
                           n2557, A => n1040, ZN => n1035);
   U628 : OAI221_X1 port map( B1 => n1947, B2 => n2525, C1 => n1944, C2 => 
                           n2493, A => n1039, ZN => n1036);
   U629 : NOR4_X1 port map( A1 => n1051, A2 => n1052, A3 => n1053, A4 => n1054,
                           ZN => n1050);
   U630 : OAI221_X1 port map( B1 => n1923, B2 => n2652, C1 => n1920, C2 => 
                           n2620, A => n1058, ZN => n1051);
   U631 : OAI221_X1 port map( B1 => n1935, B2 => n2588, C1 => n1932, C2 => 
                           n2556, A => n1057, ZN => n1052);
   U632 : OAI221_X1 port map( B1 => n1947, B2 => n2524, C1 => n1944, C2 => 
                           n2492, A => n1056, ZN => n1053);
   U633 : NOR4_X1 port map( A1 => n1068, A2 => n1069, A3 => n1070, A4 => n1071,
                           ZN => n1067);
   U634 : OAI221_X1 port map( B1 => n1923, B2 => n2651, C1 => n1920, C2 => 
                           n2619, A => n1075, ZN => n1068);
   U635 : OAI221_X1 port map( B1 => n1935, B2 => n2587, C1 => n1932, C2 => 
                           n2555, A => n1074, ZN => n1069);
   U636 : OAI221_X1 port map( B1 => n1947, B2 => n2523, C1 => n1944, C2 => 
                           n2491, A => n1073, ZN => n1070);
   U637 : NOR4_X1 port map( A1 => n1085, A2 => n1086, A3 => n1087, A4 => n1088,
                           ZN => n1084);
   U638 : OAI221_X1 port map( B1 => n1923, B2 => n2650, C1 => n1920, C2 => 
                           n2618, A => n1092, ZN => n1085);
   U639 : OAI221_X1 port map( B1 => n1935, B2 => n2586, C1 => n1932, C2 => 
                           n2554, A => n1091, ZN => n1086);
   U640 : OAI221_X1 port map( B1 => n1947, B2 => n2522, C1 => n1944, C2 => 
                           n2490, A => n1090, ZN => n1087);
   U641 : NOR4_X1 port map( A1 => n1102, A2 => n1103, A3 => n1104, A4 => n1105,
                           ZN => n1101);
   U642 : OAI221_X1 port map( B1 => n1923, B2 => n2649, C1 => n1920, C2 => 
                           n2617, A => n1117, ZN => n1102);
   U643 : OAI221_X1 port map( B1 => n1935, B2 => n2585, C1 => n1932, C2 => 
                           n2553, A => n1114, ZN => n1103);
   U644 : OAI221_X1 port map( B1 => n1947, B2 => n2521, C1 => n1944, C2 => 
                           n2489, A => n1111, ZN => n1104);
   U645 : OAI22_X1 port map( A1 => n1886, A2 => n2392, B1 => n1883, B2 => n2296
                           , ZN => n580);
   U646 : OAI22_X1 port map( A1 => n1874, A2 => n2328, B1 => n1871, B2 => n2424
                           , ZN => n585);
   U647 : OAI22_X1 port map( A1 => n1886, A2 => n2391, B1 => n1883, B2 => n2295
                           , ZN => n603);
   U648 : OAI22_X1 port map( A1 => n1874, A2 => n2327, B1 => n1871, B2 => n2423
                           , ZN => n604);
   U649 : OAI22_X1 port map( A1 => n1886, A2 => n2390, B1 => n1883, B2 => n2294
                           , ZN => n620);
   U650 : OAI22_X1 port map( A1 => n1874, A2 => n2326, B1 => n1871, B2 => n2422
                           , ZN => n621);
   U651 : OAI22_X1 port map( A1 => n1886, A2 => n2389, B1 => n1883, B2 => n2293
                           , ZN => n637);
   U652 : OAI22_X1 port map( A1 => n1874, A2 => n2325, B1 => n1871, B2 => n2421
                           , ZN => n638);
   U653 : OAI22_X1 port map( A1 => n1886, A2 => n2388, B1 => n1883, B2 => n2292
                           , ZN => n654);
   U654 : OAI22_X1 port map( A1 => n1874, A2 => n2324, B1 => n1871, B2 => n2420
                           , ZN => n655);
   U655 : OAI22_X1 port map( A1 => n1886, A2 => n2387, B1 => n1883, B2 => n2291
                           , ZN => n671);
   U656 : OAI22_X1 port map( A1 => n1874, A2 => n2323, B1 => n1871, B2 => n2419
                           , ZN => n672);
   U657 : OAI22_X1 port map( A1 => n1886, A2 => n2386, B1 => n1883, B2 => n2290
                           , ZN => n688);
   U658 : OAI22_X1 port map( A1 => n1874, A2 => n2322, B1 => n1871, B2 => n2418
                           , ZN => n689);
   U659 : OAI22_X1 port map( A1 => n1886, A2 => n2385, B1 => n1883, B2 => n2289
                           , ZN => n705);
   U660 : OAI22_X1 port map( A1 => n1874, A2 => n2321, B1 => n1871, B2 => n2417
                           , ZN => n706);
   U661 : OAI22_X1 port map( A1 => n1910, A2 => n2360, B1 => n1907, B2 => n2232
                           , ZN => n570);
   U662 : OAI22_X1 port map( A1 => n1910, A2 => n2359, B1 => n1907, B2 => n2231
                           , ZN => n601);
   U663 : OAI22_X1 port map( A1 => n1910, A2 => n2358, B1 => n1907, B2 => n2230
                           , ZN => n618);
   U664 : OAI22_X1 port map( A1 => n1910, A2 => n2357, B1 => n1907, B2 => n2229
                           , ZN => n635);
   U665 : OAI22_X1 port map( A1 => n1910, A2 => n2356, B1 => n1907, B2 => n2228
                           , ZN => n652);
   U666 : OAI22_X1 port map( A1 => n1910, A2 => n2355, B1 => n1907, B2 => n2227
                           , ZN => n669);
   U667 : OAI22_X1 port map( A1 => n1910, A2 => n2354, B1 => n1907, B2 => n2226
                           , ZN => n686);
   U668 : OAI22_X1 port map( A1 => n1910, A2 => n2353, B1 => n1907, B2 => n2225
                           , ZN => n703);
   U669 : OAI22_X1 port map( A1 => n2392, A2 => n1793, B1 => n2296, B2 => n1790
                           , ZN => n1167);
   U670 : OAI22_X1 port map( A1 => n2328, A2 => n1781, B1 => n2424, B2 => n1778
                           , ZN => n1172);
   U671 : OAI22_X1 port map( A1 => n2391, A2 => n1793, B1 => n2295, B2 => n1790
                           , ZN => n1190);
   U672 : OAI22_X1 port map( A1 => n2327, A2 => n1781, B1 => n2423, B2 => n1778
                           , ZN => n1191);
   U673 : OAI22_X1 port map( A1 => n2390, A2 => n1793, B1 => n2294, B2 => n1790
                           , ZN => n1207);
   U674 : OAI22_X1 port map( A1 => n2326, A2 => n1781, B1 => n2422, B2 => n1778
                           , ZN => n1208);
   U675 : OAI22_X1 port map( A1 => n2389, A2 => n1793, B1 => n2293, B2 => n1790
                           , ZN => n1224);
   U676 : OAI22_X1 port map( A1 => n2325, A2 => n1781, B1 => n2421, B2 => n1778
                           , ZN => n1225);
   U677 : OAI22_X1 port map( A1 => n2388, A2 => n1793, B1 => n2292, B2 => n1790
                           , ZN => n1241);
   U678 : OAI22_X1 port map( A1 => n2324, A2 => n1781, B1 => n2420, B2 => n1778
                           , ZN => n1242);
   U679 : OAI22_X1 port map( A1 => n2387, A2 => n1793, B1 => n2291, B2 => n1790
                           , ZN => n1258);
   U680 : OAI22_X1 port map( A1 => n2323, A2 => n1781, B1 => n2419, B2 => n1778
                           , ZN => n1259);
   U681 : OAI22_X1 port map( A1 => n2386, A2 => n1793, B1 => n2290, B2 => n1790
                           , ZN => n1275);
   U682 : OAI22_X1 port map( A1 => n2322, A2 => n1781, B1 => n2418, B2 => n1778
                           , ZN => n1276);
   U683 : OAI22_X1 port map( A1 => n2385, A2 => n1793, B1 => n2289, B2 => n1790
                           , ZN => n1292);
   U684 : OAI22_X1 port map( A1 => n2321, A2 => n1781, B1 => n2417, B2 => n1778
                           , ZN => n1293);
   U685 : OAI22_X1 port map( A1 => n2360, A2 => n1817, B1 => n2232, B2 => n1814
                           , ZN => n1157);
   U686 : OAI22_X1 port map( A1 => n2359, A2 => n1817, B1 => n2231, B2 => n1814
                           , ZN => n1188);
   U687 : OAI22_X1 port map( A1 => n2358, A2 => n1817, B1 => n2230, B2 => n1814
                           , ZN => n1205);
   U688 : OAI22_X1 port map( A1 => n2357, A2 => n1817, B1 => n2229, B2 => n1814
                           , ZN => n1222);
   U689 : OAI22_X1 port map( A1 => n2356, A2 => n1817, B1 => n2228, B2 => n1814
                           , ZN => n1239);
   U690 : OAI22_X1 port map( A1 => n2355, A2 => n1817, B1 => n2227, B2 => n1814
                           , ZN => n1256);
   U691 : OAI22_X1 port map( A1 => n2354, A2 => n1817, B1 => n2226, B2 => n1814
                           , ZN => n1273);
   U692 : OAI22_X1 port map( A1 => n2353, A2 => n1817, B1 => n2225, B2 => n1814
                           , ZN => n1290);
   U693 : OAI22_X1 port map( A1 => n2384, A2 => n1792, B1 => n2288, B2 => n1789
                           , ZN => n1309);
   U694 : OAI22_X1 port map( A1 => n2320, A2 => n1780, B1 => n2416, B2 => n1777
                           , ZN => n1310);
   U695 : OAI22_X1 port map( A1 => n2383, A2 => n1792, B1 => n2287, B2 => n1789
                           , ZN => n1326);
   U696 : OAI22_X1 port map( A1 => n2319, A2 => n1780, B1 => n2415, B2 => n1777
                           , ZN => n1327);
   U697 : OAI22_X1 port map( A1 => n2382, A2 => n1792, B1 => n2286, B2 => n1789
                           , ZN => n1343);
   U698 : OAI22_X1 port map( A1 => n2318, A2 => n1780, B1 => n2414, B2 => n1777
                           , ZN => n1344);
   U699 : OAI22_X1 port map( A1 => n2381, A2 => n1792, B1 => n2285, B2 => n1789
                           , ZN => n1360);
   U700 : OAI22_X1 port map( A1 => n2317, A2 => n1780, B1 => n2413, B2 => n1777
                           , ZN => n1361);
   U701 : OAI22_X1 port map( A1 => n2380, A2 => n1792, B1 => n2284, B2 => n1789
                           , ZN => n1377);
   U702 : OAI22_X1 port map( A1 => n2316, A2 => n1780, B1 => n2412, B2 => n1777
                           , ZN => n1378);
   U703 : OAI22_X1 port map( A1 => n2379, A2 => n1792, B1 => n2283, B2 => n1789
                           , ZN => n1394);
   U704 : OAI22_X1 port map( A1 => n2315, A2 => n1780, B1 => n2411, B2 => n1777
                           , ZN => n1395);
   U705 : OAI22_X1 port map( A1 => n2378, A2 => n1792, B1 => n2282, B2 => n1789
                           , ZN => n1411);
   U706 : OAI22_X1 port map( A1 => n2314, A2 => n1780, B1 => n2410, B2 => n1777
                           , ZN => n1412);
   U707 : OAI22_X1 port map( A1 => n2377, A2 => n1792, B1 => n2281, B2 => n1789
                           , ZN => n1428);
   U708 : OAI22_X1 port map( A1 => n2313, A2 => n1780, B1 => n2409, B2 => n1777
                           , ZN => n1429);
   U709 : OAI22_X1 port map( A1 => n2376, A2 => n1792, B1 => n2280, B2 => n1789
                           , ZN => n1445);
   U710 : OAI22_X1 port map( A1 => n2312, A2 => n1780, B1 => n2408, B2 => n1777
                           , ZN => n1446);
   U711 : OAI22_X1 port map( A1 => n2375, A2 => n1792, B1 => n2279, B2 => n1789
                           , ZN => n1462);
   U712 : OAI22_X1 port map( A1 => n2311, A2 => n1780, B1 => n2407, B2 => n1777
                           , ZN => n1463);
   U713 : OAI22_X1 port map( A1 => n2374, A2 => n1792, B1 => n2278, B2 => n1789
                           , ZN => n1479);
   U714 : OAI22_X1 port map( A1 => n2310, A2 => n1780, B1 => n2406, B2 => n1777
                           , ZN => n1480);
   U715 : OAI22_X1 port map( A1 => n2373, A2 => n1792, B1 => n2277, B2 => n1789
                           , ZN => n1496);
   U716 : OAI22_X1 port map( A1 => n2309, A2 => n1780, B1 => n2405, B2 => n1777
                           , ZN => n1497);
   U717 : OAI22_X1 port map( A1 => n2372, A2 => n1791, B1 => n2276, B2 => n1788
                           , ZN => n1513);
   U718 : OAI22_X1 port map( A1 => n2308, A2 => n1779, B1 => n2404, B2 => n1776
                           , ZN => n1514);
   U719 : OAI22_X1 port map( A1 => n2371, A2 => n1791, B1 => n2275, B2 => n1788
                           , ZN => n1530);
   U720 : OAI22_X1 port map( A1 => n2307, A2 => n1779, B1 => n2403, B2 => n1776
                           , ZN => n1531);
   U721 : OAI22_X1 port map( A1 => n2370, A2 => n1791, B1 => n2274, B2 => n1788
                           , ZN => n1547);
   U722 : OAI22_X1 port map( A1 => n2306, A2 => n1779, B1 => n2402, B2 => n1776
                           , ZN => n1548);
   U723 : OAI22_X1 port map( A1 => n2369, A2 => n1791, B1 => n2273, B2 => n1788
                           , ZN => n1564);
   U724 : OAI22_X1 port map( A1 => n2305, A2 => n1779, B1 => n2401, B2 => n1776
                           , ZN => n1565);
   U725 : OAI22_X1 port map( A1 => n2368, A2 => n1791, B1 => n2272, B2 => n1788
                           , ZN => n1581);
   U726 : OAI22_X1 port map( A1 => n2304, A2 => n1779, B1 => n2400, B2 => n1776
                           , ZN => n1582);
   U727 : OAI22_X1 port map( A1 => n2367, A2 => n1791, B1 => n2271, B2 => n1788
                           , ZN => n1598);
   U728 : OAI22_X1 port map( A1 => n2303, A2 => n1779, B1 => n2399, B2 => n1776
                           , ZN => n1599);
   U729 : OAI22_X1 port map( A1 => n2366, A2 => n1791, B1 => n2270, B2 => n1788
                           , ZN => n1615);
   U730 : OAI22_X1 port map( A1 => n2302, A2 => n1779, B1 => n2398, B2 => n1776
                           , ZN => n1616);
   U731 : OAI22_X1 port map( A1 => n2365, A2 => n1791, B1 => n2269, B2 => n1788
                           , ZN => n1632);
   U732 : OAI22_X1 port map( A1 => n2301, A2 => n1779, B1 => n2397, B2 => n1776
                           , ZN => n1633);
   U733 : OAI22_X1 port map( A1 => n2364, A2 => n1791, B1 => n2268, B2 => n1788
                           , ZN => n1649);
   U734 : OAI22_X1 port map( A1 => n2300, A2 => n1779, B1 => n2396, B2 => n1776
                           , ZN => n1650);
   U735 : OAI22_X1 port map( A1 => n2363, A2 => n1791, B1 => n2267, B2 => n1788
                           , ZN => n1666);
   U736 : OAI22_X1 port map( A1 => n2299, A2 => n1779, B1 => n2395, B2 => n1776
                           , ZN => n1667);
   U737 : OAI22_X1 port map( A1 => n2362, A2 => n1791, B1 => n2266, B2 => n1788
                           , ZN => n1683);
   U738 : OAI22_X1 port map( A1 => n2298, A2 => n1779, B1 => n2394, B2 => n1776
                           , ZN => n1684);
   U739 : OAI22_X1 port map( A1 => n2361, A2 => n1791, B1 => n2265, B2 => n1788
                           , ZN => n1711);
   U740 : OAI22_X1 port map( A1 => n2297, A2 => n1779, B1 => n2393, B2 => n1776
                           , ZN => n1713);
   U741 : OAI22_X1 port map( A1 => n1885, A2 => n2384, B1 => n1882, B2 => n2288
                           , ZN => n722);
   U742 : OAI22_X1 port map( A1 => n1873, A2 => n2320, B1 => n1870, B2 => n2416
                           , ZN => n723);
   U743 : OAI22_X1 port map( A1 => n1885, A2 => n2383, B1 => n1882, B2 => n2287
                           , ZN => n739);
   U744 : OAI22_X1 port map( A1 => n1873, A2 => n2319, B1 => n1870, B2 => n2415
                           , ZN => n740);
   U745 : OAI22_X1 port map( A1 => n1885, A2 => n2382, B1 => n1882, B2 => n2286
                           , ZN => n756);
   U746 : OAI22_X1 port map( A1 => n1873, A2 => n2318, B1 => n1870, B2 => n2414
                           , ZN => n757);
   U747 : OAI22_X1 port map( A1 => n1885, A2 => n2381, B1 => n1882, B2 => n2285
                           , ZN => n773);
   U748 : OAI22_X1 port map( A1 => n1873, A2 => n2317, B1 => n1870, B2 => n2413
                           , ZN => n774);
   U749 : OAI22_X1 port map( A1 => n1885, A2 => n2380, B1 => n1882, B2 => n2284
                           , ZN => n790);
   U750 : OAI22_X1 port map( A1 => n1873, A2 => n2316, B1 => n1870, B2 => n2412
                           , ZN => n791);
   U751 : OAI22_X1 port map( A1 => n1885, A2 => n2379, B1 => n1882, B2 => n2283
                           , ZN => n807);
   U752 : OAI22_X1 port map( A1 => n1873, A2 => n2315, B1 => n1870, B2 => n2411
                           , ZN => n808);
   U753 : OAI22_X1 port map( A1 => n1885, A2 => n2378, B1 => n1882, B2 => n2282
                           , ZN => n824);
   U754 : OAI22_X1 port map( A1 => n1873, A2 => n2314, B1 => n1870, B2 => n2410
                           , ZN => n825);
   U755 : OAI22_X1 port map( A1 => n1885, A2 => n2377, B1 => n1882, B2 => n2281
                           , ZN => n841);
   U756 : OAI22_X1 port map( A1 => n1873, A2 => n2313, B1 => n1870, B2 => n2409
                           , ZN => n842);
   U757 : OAI22_X1 port map( A1 => n1885, A2 => n2376, B1 => n1882, B2 => n2280
                           , ZN => n858);
   U758 : OAI22_X1 port map( A1 => n1873, A2 => n2312, B1 => n1870, B2 => n2408
                           , ZN => n859);
   U759 : OAI22_X1 port map( A1 => n1885, A2 => n2375, B1 => n1882, B2 => n2279
                           , ZN => n875);
   U760 : OAI22_X1 port map( A1 => n1873, A2 => n2311, B1 => n1870, B2 => n2407
                           , ZN => n876);
   U761 : OAI22_X1 port map( A1 => n1885, A2 => n2374, B1 => n1882, B2 => n2278
                           , ZN => n892);
   U762 : OAI22_X1 port map( A1 => n1873, A2 => n2310, B1 => n1870, B2 => n2406
                           , ZN => n893);
   U763 : OAI22_X1 port map( A1 => n1885, A2 => n2373, B1 => n1882, B2 => n2277
                           , ZN => n909);
   U764 : OAI22_X1 port map( A1 => n1873, A2 => n2309, B1 => n1870, B2 => n2405
                           , ZN => n910);
   U765 : OAI22_X1 port map( A1 => n1884, A2 => n2372, B1 => n1881, B2 => n2276
                           , ZN => n926);
   U766 : OAI22_X1 port map( A1 => n1872, A2 => n2308, B1 => n1869, B2 => n2404
                           , ZN => n927);
   U767 : OAI22_X1 port map( A1 => n1884, A2 => n2371, B1 => n1881, B2 => n2275
                           , ZN => n943);
   U768 : OAI22_X1 port map( A1 => n1872, A2 => n2307, B1 => n1869, B2 => n2403
                           , ZN => n944);
   U769 : OAI22_X1 port map( A1 => n1884, A2 => n2370, B1 => n1881, B2 => n2274
                           , ZN => n960);
   U770 : OAI22_X1 port map( A1 => n1872, A2 => n2306, B1 => n1869, B2 => n2402
                           , ZN => n961);
   U771 : OAI22_X1 port map( A1 => n1884, A2 => n2369, B1 => n1881, B2 => n2273
                           , ZN => n977);
   U772 : OAI22_X1 port map( A1 => n1872, A2 => n2305, B1 => n1869, B2 => n2401
                           , ZN => n978);
   U773 : OAI22_X1 port map( A1 => n1884, A2 => n2368, B1 => n1881, B2 => n2272
                           , ZN => n994);
   U774 : OAI22_X1 port map( A1 => n1872, A2 => n2304, B1 => n1869, B2 => n2400
                           , ZN => n995);
   U775 : OAI22_X1 port map( A1 => n1884, A2 => n2367, B1 => n1881, B2 => n2271
                           , ZN => n1011);
   U776 : OAI22_X1 port map( A1 => n1872, A2 => n2303, B1 => n1869, B2 => n2399
                           , ZN => n1012);
   U777 : OAI22_X1 port map( A1 => n1884, A2 => n2366, B1 => n1881, B2 => n2270
                           , ZN => n1028);
   U778 : OAI22_X1 port map( A1 => n1872, A2 => n2302, B1 => n1869, B2 => n2398
                           , ZN => n1029);
   U779 : OAI22_X1 port map( A1 => n1884, A2 => n2365, B1 => n1881, B2 => n2269
                           , ZN => n1045);
   U780 : OAI22_X1 port map( A1 => n1872, A2 => n2301, B1 => n1869, B2 => n2397
                           , ZN => n1046);
   U781 : OAI22_X1 port map( A1 => n1884, A2 => n2364, B1 => n1881, B2 => n2268
                           , ZN => n1062);
   U782 : OAI22_X1 port map( A1 => n1872, A2 => n2300, B1 => n1869, B2 => n2396
                           , ZN => n1063);
   U783 : OAI22_X1 port map( A1 => n1884, A2 => n2363, B1 => n1881, B2 => n2267
                           , ZN => n1079);
   U784 : OAI22_X1 port map( A1 => n1872, A2 => n2299, B1 => n1869, B2 => n2395
                           , ZN => n1080);
   U785 : OAI22_X1 port map( A1 => n1884, A2 => n2362, B1 => n1881, B2 => n2266
                           , ZN => n1096);
   U786 : OAI22_X1 port map( A1 => n1872, A2 => n2298, B1 => n1869, B2 => n2394
                           , ZN => n1097);
   U787 : OAI22_X1 port map( A1 => n1884, A2 => n2361, B1 => n1881, B2 => n2265
                           , ZN => n1124);
   U788 : OAI22_X1 port map( A1 => n1872, A2 => n2297, B1 => n1869, B2 => n2393
                           , ZN => n1126);
   U789 : OAI22_X1 port map( A1 => n2352, A2 => n1816, B1 => n2224, B2 => n1813
                           , ZN => n1307);
   U790 : OAI22_X1 port map( A1 => n2351, A2 => n1816, B1 => n2223, B2 => n1813
                           , ZN => n1324);
   U791 : OAI22_X1 port map( A1 => n2350, A2 => n1816, B1 => n2222, B2 => n1813
                           , ZN => n1341);
   U792 : OAI22_X1 port map( A1 => n2349, A2 => n1816, B1 => n2221, B2 => n1813
                           , ZN => n1358);
   U793 : OAI22_X1 port map( A1 => n2348, A2 => n1816, B1 => n2220, B2 => n1813
                           , ZN => n1375);
   U794 : OAI22_X1 port map( A1 => n2347, A2 => n1816, B1 => n2219, B2 => n1813
                           , ZN => n1392);
   U795 : OAI22_X1 port map( A1 => n2346, A2 => n1816, B1 => n2218, B2 => n1813
                           , ZN => n1409);
   U796 : OAI22_X1 port map( A1 => n2345, A2 => n1816, B1 => n2217, B2 => n1813
                           , ZN => n1426);
   U797 : OAI22_X1 port map( A1 => n2344, A2 => n1816, B1 => n2216, B2 => n1813
                           , ZN => n1443);
   U798 : OAI22_X1 port map( A1 => n2343, A2 => n1816, B1 => n2215, B2 => n1813
                           , ZN => n1460);
   U799 : OAI22_X1 port map( A1 => n2342, A2 => n1816, B1 => n2214, B2 => n1813
                           , ZN => n1477);
   U800 : OAI22_X1 port map( A1 => n2341, A2 => n1816, B1 => n2213, B2 => n1813
                           , ZN => n1494);
   U801 : OAI22_X1 port map( A1 => n2340, A2 => n1815, B1 => n2212, B2 => n1812
                           , ZN => n1511);
   U802 : OAI22_X1 port map( A1 => n2339, A2 => n1815, B1 => n2211, B2 => n1812
                           , ZN => n1528);
   U803 : OAI22_X1 port map( A1 => n2338, A2 => n1815, B1 => n2210, B2 => n1812
                           , ZN => n1545);
   U804 : OAI22_X1 port map( A1 => n2337, A2 => n1815, B1 => n2209, B2 => n1812
                           , ZN => n1562);
   U805 : OAI22_X1 port map( A1 => n2336, A2 => n1815, B1 => n2208, B2 => n1812
                           , ZN => n1579);
   U806 : OAI22_X1 port map( A1 => n2335, A2 => n1815, B1 => n2207, B2 => n1812
                           , ZN => n1596);
   U807 : OAI22_X1 port map( A1 => n2334, A2 => n1815, B1 => n2206, B2 => n1812
                           , ZN => n1613);
   U808 : OAI22_X1 port map( A1 => n2333, A2 => n1815, B1 => n2205, B2 => n1812
                           , ZN => n1630);
   U809 : OAI22_X1 port map( A1 => n2332, A2 => n1815, B1 => n2204, B2 => n1812
                           , ZN => n1647);
   U810 : OAI22_X1 port map( A1 => n2331, A2 => n1815, B1 => n2203, B2 => n1812
                           , ZN => n1664);
   U811 : OAI22_X1 port map( A1 => n2330, A2 => n1815, B1 => n2202, B2 => n1812
                           , ZN => n1681);
   U812 : OAI22_X1 port map( A1 => n2329, A2 => n1815, B1 => n2201, B2 => n1812
                           , ZN => n1706);
   U813 : OAI22_X1 port map( A1 => n1909, A2 => n2352, B1 => n1906, B2 => n2224
                           , ZN => n720);
   U814 : OAI22_X1 port map( A1 => n1909, A2 => n2351, B1 => n1906, B2 => n2223
                           , ZN => n737);
   U815 : OAI22_X1 port map( A1 => n1909, A2 => n2350, B1 => n1906, B2 => n2222
                           , ZN => n754);
   U816 : OAI22_X1 port map( A1 => n1909, A2 => n2349, B1 => n1906, B2 => n2221
                           , ZN => n771);
   U817 : OAI22_X1 port map( A1 => n1909, A2 => n2348, B1 => n1906, B2 => n2220
                           , ZN => n788);
   U818 : OAI22_X1 port map( A1 => n1909, A2 => n2347, B1 => n1906, B2 => n2219
                           , ZN => n805);
   U819 : OAI22_X1 port map( A1 => n1909, A2 => n2346, B1 => n1906, B2 => n2218
                           , ZN => n822);
   U820 : OAI22_X1 port map( A1 => n1909, A2 => n2345, B1 => n1906, B2 => n2217
                           , ZN => n839);
   U821 : OAI22_X1 port map( A1 => n1909, A2 => n2344, B1 => n1906, B2 => n2216
                           , ZN => n856);
   U822 : OAI22_X1 port map( A1 => n1909, A2 => n2343, B1 => n1906, B2 => n2215
                           , ZN => n873);
   U823 : OAI22_X1 port map( A1 => n1909, A2 => n2342, B1 => n1906, B2 => n2214
                           , ZN => n890);
   U824 : OAI22_X1 port map( A1 => n1909, A2 => n2341, B1 => n1906, B2 => n2213
                           , ZN => n907);
   U825 : OAI22_X1 port map( A1 => n1908, A2 => n2340, B1 => n1905, B2 => n2212
                           , ZN => n924);
   U826 : OAI22_X1 port map( A1 => n1908, A2 => n2339, B1 => n1905, B2 => n2211
                           , ZN => n941);
   U827 : OAI22_X1 port map( A1 => n1908, A2 => n2338, B1 => n1905, B2 => n2210
                           , ZN => n958);
   U828 : OAI22_X1 port map( A1 => n1908, A2 => n2337, B1 => n1905, B2 => n2209
                           , ZN => n975);
   U829 : OAI22_X1 port map( A1 => n1908, A2 => n2336, B1 => n1905, B2 => n2208
                           , ZN => n992);
   U830 : OAI22_X1 port map( A1 => n1908, A2 => n2335, B1 => n1905, B2 => n2207
                           , ZN => n1009);
   U831 : OAI22_X1 port map( A1 => n1908, A2 => n2334, B1 => n1905, B2 => n2206
                           , ZN => n1026);
   U832 : OAI22_X1 port map( A1 => n1908, A2 => n2333, B1 => n1905, B2 => n2205
                           , ZN => n1043);
   U833 : OAI22_X1 port map( A1 => n1908, A2 => n2332, B1 => n1905, B2 => n2204
                           , ZN => n1060);
   U834 : OAI22_X1 port map( A1 => n1908, A2 => n2331, B1 => n1905, B2 => n2203
                           , ZN => n1077);
   U835 : OAI22_X1 port map( A1 => n1908, A2 => n2330, B1 => n1905, B2 => n2202
                           , ZN => n1094);
   U836 : OAI22_X1 port map( A1 => n1908, A2 => n2329, B1 => n1905, B2 => n2201
                           , ZN => n1119);
   U837 : NAND2_X1 port map( A1 => n1697, A2 => n1702, ZN => n1146);
   U838 : NAND2_X1 port map( A1 => n1697, A2 => n1703, ZN => n1145);
   U839 : NAND2_X1 port map( A1 => n1110, A2 => n1116, ZN => n558);
   U840 : NAND2_X1 port map( A1 => n1110, A2 => n1115, ZN => n559);
   U841 : NAND2_X1 port map( A1 => n1700, A2 => n1703, ZN => n1150);
   U842 : NAND2_X1 port map( A1 => n1113, A2 => n1116, ZN => n563);
   U843 : NAND2_X1 port map( A1 => n1708, A2 => n1695, ZN => n1169);
   U844 : NAND2_X1 port map( A1 => n1708, A2 => n1699, ZN => n1174);
   U845 : NAND2_X1 port map( A1 => n1708, A2 => n1697, ZN => n1158);
   U846 : NAND2_X1 port map( A1 => n1121, A2 => n1108, ZN => n582);
   U847 : NAND2_X1 port map( A1 => n1121, A2 => n1112, ZN => n587);
   U848 : NAND2_X1 port map( A1 => n1121, A2 => n1110, ZN => n571);
   U849 : NAND2_X1 port map( A1 => n1712, A2 => n1697, ZN => n1168);
   U850 : NAND2_X1 port map( A1 => n1712, A2 => n1695, ZN => n1173);
   U851 : NAND2_X1 port map( A1 => n1710, A2 => n1699, ZN => n1161);
   U852 : NAND2_X1 port map( A1 => n1710, A2 => n1695, ZN => n1160);
   U853 : NAND2_X1 port map( A1 => n1125, A2 => n1110, ZN => n581);
   U854 : NAND2_X1 port map( A1 => n1125, A2 => n1108, ZN => n586);
   U855 : NAND2_X1 port map( A1 => n1123, A2 => n1108, ZN => n573);
   U856 : NAND2_X1 port map( A1 => n1123, A2 => n1112, ZN => n574);
   U857 : NAND2_X1 port map( A1 => n1694, A2 => n1697, ZN => n1136);
   U858 : NAND2_X1 port map( A1 => n1696, A2 => n1697, ZN => n1135);
   U859 : NAND2_X1 port map( A1 => n1109, A2 => n1110, ZN => n548);
   U860 : NAND2_X1 port map( A1 => n1107, A2 => n1110, ZN => n549);
   U861 : NAND2_X1 port map( A1 => n1707, A2 => n1700, ZN => n1159);
   U862 : NAND2_X1 port map( A1 => n1694, A2 => n1700, ZN => n1141);
   U863 : NAND2_X1 port map( A1 => n1696, A2 => n1700, ZN => n1140);
   U864 : NAND2_X1 port map( A1 => n1702, A2 => n1700, ZN => n1151);
   U865 : NAND2_X1 port map( A1 => n1109, A2 => n1113, ZN => n553);
   U866 : NAND2_X1 port map( A1 => n1107, A2 => n1113, ZN => n554);
   U867 : NAND2_X1 port map( A1 => n1115, A2 => n1113, ZN => n564);
   U868 : NAND2_X1 port map( A1 => n1120, A2 => n1113, ZN => n572);
   U869 : AND2_X1 port map( A1 => n1708, A2 => n1700, ZN => n1166);
   U870 : AND2_X1 port map( A1 => n1121, A2 => n1113, ZN => n579);
   U871 : AND2_X1 port map( A1 => n1699, A2 => n1703, ZN => n1153);
   U872 : AND2_X1 port map( A1 => n1699, A2 => n1702, ZN => n1154);
   U873 : AND2_X1 port map( A1 => n1112, A2 => n1116, ZN => n566);
   U874 : AND2_X1 port map( A1 => n1112, A2 => n1115, ZN => n567);
   U875 : AND2_X1 port map( A1 => n1710, A2 => n1697, ZN => n1163);
   U876 : AND2_X1 port map( A1 => n1712, A2 => n1699, ZN => n1165);
   U877 : AND2_X1 port map( A1 => n1712, A2 => n1700, ZN => n1170);
   U878 : AND2_X1 port map( A1 => n1710, A2 => n1700, ZN => n1155);
   U879 : AND2_X1 port map( A1 => n1108, A2 => n1116, ZN => n561);
   U880 : AND2_X1 port map( A1 => n1108, A2 => n1115, ZN => n562);
   U881 : AND2_X1 port map( A1 => n1695, A2 => n1703, ZN => n1148);
   U882 : AND2_X1 port map( A1 => n1695, A2 => n1702, ZN => n1149);
   U883 : AND2_X1 port map( A1 => n1123, A2 => n1110, ZN => n576);
   U884 : AND2_X1 port map( A1 => n1707, A2 => n1697, ZN => n1171);
   U885 : AND2_X1 port map( A1 => n1120, A2 => n1110, ZN => n584);
   U886 : AND2_X1 port map( A1 => n1125, A2 => n1112, ZN => n578);
   U887 : AND2_X1 port map( A1 => n1125, A2 => n1113, ZN => n583);
   U888 : AND2_X1 port map( A1 => n1123, A2 => n1113, ZN => n568);
   U889 : AND2_X1 port map( A1 => n1696, A2 => n1699, ZN => n1143);
   U890 : AND2_X1 port map( A1 => n1694, A2 => n1699, ZN => n1144);
   U891 : AND2_X1 port map( A1 => n1707, A2 => n1699, ZN => n1164);
   U892 : AND2_X1 port map( A1 => n1109, A2 => n1112, ZN => n556);
   U893 : AND2_X1 port map( A1 => n1107, A2 => n1112, ZN => n557);
   U894 : AND2_X1 port map( A1 => n1120, A2 => n1112, ZN => n577);
   U895 : AND2_X1 port map( A1 => n1109, A2 => n1108, ZN => n551);
   U896 : AND2_X1 port map( A1 => n1107, A2 => n1108, ZN => n552);
   U897 : AND2_X1 port map( A1 => n1696, A2 => n1695, ZN => n1138);
   U898 : AND2_X1 port map( A1 => n1694, A2 => n1695, ZN => n1139);
   U899 : OAI21_X1 port map( B1 => n533, B2 => n539, A => n2161, ZN => N340);
   U900 : OAI21_X1 port map( B1 => n532, B2 => n539, A => n2161, ZN => N341);
   U901 : OAI21_X1 port map( B1 => n531, B2 => n539, A => n2161, ZN => N342);
   U902 : OAI21_X1 port map( B1 => n530, B2 => n539, A => n2161, ZN => N343);
   U903 : OAI21_X1 port map( B1 => n529, B2 => n539, A => n2161, ZN => N344);
   U904 : OAI21_X1 port map( B1 => n528, B2 => n539, A => n2161, ZN => N345);
   U905 : OAI21_X1 port map( B1 => n534, B2 => n538, A => n2161, ZN => N347);
   U906 : OAI21_X1 port map( B1 => n534, B2 => n539, A => n2159, ZN => N307);
   U907 : OAI21_X1 port map( B1 => n537, B2 => n539, A => n2160, ZN => N346);
   U908 : OAI21_X1 port map( B1 => n533, B2 => n538, A => n2160, ZN => N348);
   U909 : OAI21_X1 port map( B1 => n532, B2 => n538, A => n2160, ZN => N349);
   U910 : OAI21_X1 port map( B1 => n531, B2 => n538, A => n2160, ZN => N350);
   U911 : OAI21_X1 port map( B1 => n530, B2 => n538, A => n2160, ZN => N351);
   U912 : OAI21_X1 port map( B1 => n529, B2 => n538, A => n2160, ZN => N352);
   U913 : OAI21_X1 port map( B1 => n528, B2 => n538, A => n2160, ZN => N353);
   U914 : OAI21_X1 port map( B1 => n537, B2 => n538, A => n2160, ZN => N354);
   U915 : OAI21_X1 port map( B1 => n534, B2 => n536, A => n2160, ZN => N355);
   U916 : OAI21_X1 port map( B1 => n533, B2 => n536, A => n2160, ZN => N356);
   U917 : OAI21_X1 port map( B1 => n532, B2 => n536, A => n2160, ZN => N357);
   U918 : OAI21_X1 port map( B1 => n531, B2 => n536, A => n2159, ZN => N358);
   U919 : OAI21_X1 port map( B1 => n530, B2 => n536, A => n2160, ZN => N359);
   U920 : OAI21_X1 port map( B1 => n529, B2 => n536, A => n2159, ZN => N360);
   U921 : OAI21_X1 port map( B1 => n528, B2 => n536, A => n2159, ZN => N361);
   U922 : OAI21_X1 port map( B1 => n536, B2 => n537, A => n2159, ZN => N362);
   U923 : OAI21_X1 port map( B1 => n527, B2 => n534, A => n2159, ZN => N363);
   U924 : OAI21_X1 port map( B1 => n527, B2 => n533, A => n2159, ZN => N364);
   U925 : OAI21_X1 port map( B1 => n527, B2 => n532, A => n2159, ZN => N365);
   U926 : OAI21_X1 port map( B1 => n527, B2 => n531, A => n2159, ZN => N366);
   U927 : OAI21_X1 port map( B1 => n527, B2 => n530, A => n2159, ZN => N367);
   U928 : OAI21_X1 port map( B1 => n527, B2 => n529, A => n2159, ZN => N368);
   U929 : OAI21_X1 port map( B1 => n527, B2 => n528, A => n2159, ZN => N369);
   U930 : AND2_X1 port map( A1 => n2689, A2 => n2162, ZN => N371);
   U931 : AND2_X1 port map( A1 => datain(0), A2 => n2161, ZN => N308);
   U932 : AND2_X1 port map( A1 => datain(15), A2 => n2161, ZN => N323);
   U933 : AND2_X1 port map( A1 => datain(26), A2 => n2161, ZN => N334);
   U934 : AND2_X1 port map( A1 => datain(27), A2 => n2161, ZN => N335);
   U935 : AND2_X1 port map( A1 => datain(28), A2 => n2161, ZN => N336);
   U936 : AND2_X1 port map( A1 => datain(29), A2 => n2161, ZN => N337);
   U937 : AND2_X1 port map( A1 => datain(30), A2 => n2161, ZN => N338);
   U938 : AND2_X1 port map( A1 => datain(31), A2 => n2161, ZN => N339);
   U939 : AND2_X1 port map( A1 => datain(8), A2 => n2162, ZN => N316);
   U940 : AND2_X1 port map( A1 => datain(9), A2 => n2162, ZN => N317);
   U941 : AND2_X1 port map( A1 => datain(10), A2 => n2162, ZN => N318);
   U942 : AND2_X1 port map( A1 => datain(11), A2 => n2162, ZN => N319);
   U943 : AND2_X1 port map( A1 => datain(12), A2 => n2162, ZN => N320);
   U944 : AND2_X1 port map( A1 => datain(13), A2 => n2162, ZN => N321);
   U945 : AND2_X1 port map( A1 => datain(14), A2 => n2162, ZN => N322);
   U946 : AND2_X1 port map( A1 => datain(16), A2 => n2162, ZN => N324);
   U947 : AND2_X1 port map( A1 => datain(17), A2 => n2162, ZN => N325);
   U948 : AND2_X1 port map( A1 => datain(18), A2 => n2162, ZN => N326);
   U949 : AND2_X1 port map( A1 => datain(19), A2 => n2162, ZN => N327);
   U950 : AND2_X1 port map( A1 => datain(20), A2 => n2162, ZN => N328);
   U951 : AND2_X1 port map( A1 => datain(21), A2 => n2162, ZN => N329);
   U952 : AND2_X1 port map( A1 => datain(22), A2 => n2162, ZN => N330);
   U953 : AND2_X1 port map( A1 => datain(23), A2 => n2162, ZN => N331);
   U954 : AND2_X1 port map( A1 => datain(24), A2 => n2162, ZN => N332);
   U955 : AND2_X1 port map( A1 => datain(25), A2 => n2162, ZN => N333);
   U956 : AND2_X1 port map( A1 => datain(1), A2 => n2163, ZN => N309);
   U957 : AND2_X1 port map( A1 => datain(2), A2 => n2163, ZN => N310);
   U958 : AND2_X1 port map( A1 => datain(3), A2 => n2163, ZN => N311);
   U959 : AND2_X1 port map( A1 => datain(4), A2 => n2163, ZN => N312);
   U960 : AND2_X1 port map( A1 => datain(5), A2 => n2163, ZN => N313);
   U961 : AND2_X1 port map( A1 => datain(6), A2 => n2163, ZN => N314);
   U962 : AND2_X1 port map( A1 => datain(7), A2 => n2163, ZN => N315);
   U963 : NOR2_X1 port map( A1 => n2682, A2 => add_rd1(1), ZN => n1700);
   U964 : NOR2_X1 port map( A1 => n2686, A2 => add_rd2(1), ZN => n1113);
   U965 : NOR3_X1 port map( A1 => add_rd1(0), A2 => add_rd1(4), A3 => n2681, ZN
                           => n1708);
   U966 : NOR3_X1 port map( A1 => add_rd2(0), A2 => add_rd2(4), A3 => n2685, ZN
                           => n1121);
   U967 : NOR3_X1 port map( A1 => add_rd1(3), A2 => add_rd1(4), A3 => n2684, ZN
                           => n1710);
   U968 : NOR3_X1 port map( A1 => n2684, A2 => add_rd1(4), A3 => n2681, ZN => 
                           n1712);
   U969 : NOR2_X1 port map( A1 => add_rd2(1), A2 => add_rd2(2), ZN => n1108);
   U970 : NOR2_X1 port map( A1 => add_rd1(1), A2 => add_rd1(2), ZN => n1695);
   U971 : NOR3_X1 port map( A1 => add_rd2(3), A2 => add_rd2(4), A3 => n2688, ZN
                           => n1123);
   U972 : NOR3_X1 port map( A1 => n2688, A2 => add_rd2(4), A3 => n2685, ZN => 
                           n1125);
   U973 : NOR3_X1 port map( A1 => add_rd1(3), A2 => add_rd1(4), A3 => 
                           add_rd1(0), ZN => n1707);
   U974 : NOR3_X1 port map( A1 => add_rd2(3), A2 => add_rd2(4), A3 => 
                           add_rd2(0), ZN => n1120);
   U975 : OAI221_X1 port map( B1 => n1961, B2 => n2488, C1 => n1958, C2 => 
                           n2456, A => n550, ZN => n547);
   U976 : AOI22_X1 port map( A1 => registers_17_0_port, A2 => n1955, B1 => 
                           registers_16_0_port, B2 => n1952, ZN => n550);
   U977 : OAI221_X1 port map( B1 => n1961, B2 => n2487, C1 => n1958, C2 => 
                           n2455, A => n596, ZN => n595);
   U978 : AOI22_X1 port map( A1 => registers_17_1_port, A2 => n1955, B1 => 
                           registers_16_1_port, B2 => n1952, ZN => n596);
   U979 : OAI221_X1 port map( B1 => n1961, B2 => n2486, C1 => n1958, C2 => 
                           n2454, A => n613, ZN => n612);
   U980 : AOI22_X1 port map( A1 => registers_17_2_port, A2 => n1955, B1 => 
                           registers_16_2_port, B2 => n1952, ZN => n613);
   U981 : OAI221_X1 port map( B1 => n1961, B2 => n2485, C1 => n1958, C2 => 
                           n2453, A => n630, ZN => n629);
   U982 : AOI22_X1 port map( A1 => registers_17_3_port, A2 => n1955, B1 => 
                           registers_16_3_port, B2 => n1952, ZN => n630);
   U983 : OAI221_X1 port map( B1 => n1961, B2 => n2484, C1 => n1958, C2 => 
                           n2452, A => n647, ZN => n646);
   U984 : AOI22_X1 port map( A1 => registers_17_4_port, A2 => n1955, B1 => 
                           registers_16_4_port, B2 => n1952, ZN => n647);
   U985 : OAI221_X1 port map( B1 => n1961, B2 => n2483, C1 => n1958, C2 => 
                           n2451, A => n664, ZN => n663);
   U986 : AOI22_X1 port map( A1 => registers_17_5_port, A2 => n1955, B1 => 
                           registers_16_5_port, B2 => n1952, ZN => n664);
   U987 : OAI221_X1 port map( B1 => n1961, B2 => n2482, C1 => n1958, C2 => 
                           n2450, A => n681, ZN => n680);
   U988 : AOI22_X1 port map( A1 => registers_17_6_port, A2 => n1955, B1 => 
                           registers_16_6_port, B2 => n1952, ZN => n681);
   U989 : OAI221_X1 port map( B1 => n1961, B2 => n2481, C1 => n1958, C2 => 
                           n2449, A => n698, ZN => n697);
   U990 : AOI22_X1 port map( A1 => registers_17_7_port, A2 => n1955, B1 => 
                           registers_16_7_port, B2 => n1952, ZN => n698);
   U991 : OAI221_X1 port map( B1 => n2488, B2 => n1868, C1 => n2456, C2 => 
                           n1865, A => n1137, ZN => n1134);
   U992 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_0_port, B1 => 
                           n1857, B2 => registers_16_0_port, ZN => n1137);
   U993 : OAI221_X1 port map( B1 => n2487, B2 => n1868, C1 => n2455, C2 => 
                           n1865, A => n1183, ZN => n1182);
   U994 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_1_port, B1 => 
                           n1857, B2 => registers_16_1_port, ZN => n1183);
   U995 : OAI221_X1 port map( B1 => n2486, B2 => n1868, C1 => n2454, C2 => 
                           n1865, A => n1200, ZN => n1199);
   U996 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_2_port, B1 => 
                           n1857, B2 => registers_16_2_port, ZN => n1200);
   U997 : OAI221_X1 port map( B1 => n2485, B2 => n1868, C1 => n2453, C2 => 
                           n1865, A => n1217, ZN => n1216);
   U998 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_3_port, B1 => 
                           n1857, B2 => registers_16_3_port, ZN => n1217);
   U999 : OAI221_X1 port map( B1 => n2484, B2 => n1868, C1 => n2452, C2 => 
                           n1865, A => n1234, ZN => n1233);
   U1000 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_4_port, B1 => 
                           n1857, B2 => registers_16_4_port, ZN => n1234);
   U1001 : OAI221_X1 port map( B1 => n2483, B2 => n1868, C1 => n2451, C2 => 
                           n1865, A => n1251, ZN => n1250);
   U1002 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_5_port, B1 => 
                           n1857, B2 => registers_16_5_port, ZN => n1251);
   U1003 : OAI221_X1 port map( B1 => n2482, B2 => n1868, C1 => n2450, C2 => 
                           n1865, A => n1268, ZN => n1267);
   U1004 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_6_port, B1 => 
                           n1857, B2 => registers_16_6_port, ZN => n1268);
   U1005 : OAI221_X1 port map( B1 => n2481, B2 => n1868, C1 => n2449, C2 => 
                           n1865, A => n1285, ZN => n1284);
   U1006 : AOI22_X1 port map( A1 => n1862, A2 => registers_17_7_port, B1 => 
                           n1857, B2 => registers_16_7_port, ZN => n1285);
   U1007 : OAI221_X1 port map( B1 => n2480, B2 => n1867, C1 => n2448, C2 => 
                           n1864, A => n1302, ZN => n1301);
   U1008 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_8_port, B1 => 
                           n1857, B2 => registers_16_8_port, ZN => n1302);
   U1009 : OAI221_X1 port map( B1 => n2479, B2 => n1867, C1 => n2447, C2 => 
                           n1864, A => n1319, ZN => n1318);
   U1010 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_9_port, B1 => 
                           n1857, B2 => registers_16_9_port, ZN => n1319);
   U1011 : OAI221_X1 port map( B1 => n2478, B2 => n1867, C1 => n2446, C2 => 
                           n1864, A => n1336, ZN => n1335);
   U1012 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_10_port, B1 => 
                           n1857, B2 => registers_16_10_port, ZN => n1336);
   U1013 : OAI221_X1 port map( B1 => n2477, B2 => n1867, C1 => n2445, C2 => 
                           n1864, A => n1353, ZN => n1352);
   U1014 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_11_port, B1 => 
                           n1857, B2 => registers_16_11_port, ZN => n1353);
   U1015 : OAI221_X1 port map( B1 => n2476, B2 => n1867, C1 => n2444, C2 => 
                           n1864, A => n1370, ZN => n1369);
   U1016 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_12_port, B1 => 
                           n1858, B2 => registers_16_12_port, ZN => n1370);
   U1017 : OAI221_X1 port map( B1 => n2475, B2 => n1867, C1 => n2443, C2 => 
                           n1864, A => n1387, ZN => n1386);
   U1018 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_13_port, B1 => 
                           n1858, B2 => registers_16_13_port, ZN => n1387);
   U1019 : OAI221_X1 port map( B1 => n2474, B2 => n1867, C1 => n2442, C2 => 
                           n1864, A => n1404, ZN => n1403);
   U1020 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_14_port, B1 => 
                           n1858, B2 => registers_16_14_port, ZN => n1404);
   U1021 : OAI221_X1 port map( B1 => n2473, B2 => n1867, C1 => n2441, C2 => 
                           n1864, A => n1421, ZN => n1420);
   U1022 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_15_port, B1 => 
                           n1858, B2 => registers_16_15_port, ZN => n1421);
   U1023 : OAI221_X1 port map( B1 => n2472, B2 => n1867, C1 => n2440, C2 => 
                           n1864, A => n1438, ZN => n1437);
   U1024 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_16_port, B1 => 
                           n1858, B2 => registers_16_16_port, ZN => n1438);
   U1025 : OAI221_X1 port map( B1 => n2471, B2 => n1867, C1 => n2439, C2 => 
                           n1864, A => n1455, ZN => n1454);
   U1026 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_17_port, B1 => 
                           n1858, B2 => registers_16_17_port, ZN => n1455);
   U1027 : OAI221_X1 port map( B1 => n2470, B2 => n1867, C1 => n2438, C2 => 
                           n1864, A => n1472, ZN => n1471);
   U1028 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_18_port, B1 => 
                           n1858, B2 => registers_16_18_port, ZN => n1472);
   U1029 : OAI221_X1 port map( B1 => n2469, B2 => n1867, C1 => n2437, C2 => 
                           n1864, A => n1489, ZN => n1488);
   U1030 : AOI22_X1 port map( A1 => n1861, A2 => registers_17_19_port, B1 => 
                           n1858, B2 => registers_16_19_port, ZN => n1489);
   U1031 : OAI221_X1 port map( B1 => n2468, B2 => n1866, C1 => n2436, C2 => 
                           n1863, A => n1506, ZN => n1505);
   U1032 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_20_port, B1 => 
                           n1858, B2 => registers_16_20_port, ZN => n1506);
   U1033 : OAI221_X1 port map( B1 => n2467, B2 => n1866, C1 => n2435, C2 => 
                           n1863, A => n1523, ZN => n1522);
   U1034 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_21_port, B1 => 
                           n1858, B2 => registers_16_21_port, ZN => n1523);
   U1035 : OAI221_X1 port map( B1 => n2466, B2 => n1866, C1 => n2434, C2 => 
                           n1863, A => n1540, ZN => n1539);
   U1036 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_22_port, B1 => 
                           n1858, B2 => registers_16_22_port, ZN => n1540);
   U1037 : OAI221_X1 port map( B1 => n2465, B2 => n1866, C1 => n2433, C2 => 
                           n1863, A => n1557, ZN => n1556);
   U1038 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_23_port, B1 => 
                           n1858, B2 => registers_16_23_port, ZN => n1557);
   U1039 : OAI221_X1 port map( B1 => n2464, B2 => n1866, C1 => n2432, C2 => 
                           n1863, A => n1574, ZN => n1573);
   U1040 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_24_port, B1 => 
                           n1859, B2 => registers_16_24_port, ZN => n1574);
   U1041 : OAI221_X1 port map( B1 => n2463, B2 => n1866, C1 => n2431, C2 => 
                           n1863, A => n1591, ZN => n1590);
   U1042 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_25_port, B1 => 
                           n1859, B2 => registers_16_25_port, ZN => n1591);
   U1043 : OAI221_X1 port map( B1 => n2462, B2 => n1866, C1 => n2430, C2 => 
                           n1863, A => n1608, ZN => n1607);
   U1044 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_26_port, B1 => 
                           n1859, B2 => registers_16_26_port, ZN => n1608);
   U1045 : OAI221_X1 port map( B1 => n2461, B2 => n1866, C1 => n2429, C2 => 
                           n1863, A => n1625, ZN => n1624);
   U1046 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_27_port, B1 => 
                           n1859, B2 => registers_16_27_port, ZN => n1625);
   U1047 : OAI221_X1 port map( B1 => n2460, B2 => n1866, C1 => n2428, C2 => 
                           n1863, A => n1642, ZN => n1641);
   U1048 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_28_port, B1 => 
                           n1859, B2 => registers_16_28_port, ZN => n1642);
   U1049 : OAI221_X1 port map( B1 => n2459, B2 => n1866, C1 => n2427, C2 => 
                           n1863, A => n1659, ZN => n1658);
   U1050 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_29_port, B1 => 
                           n1859, B2 => registers_16_29_port, ZN => n1659);
   U1051 : OAI221_X1 port map( B1 => n2458, B2 => n1866, C1 => n2426, C2 => 
                           n1863, A => n1676, ZN => n1675);
   U1052 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_30_port, B1 => 
                           n1859, B2 => registers_16_30_port, ZN => n1676);
   U1053 : OAI221_X1 port map( B1 => n2457, B2 => n1866, C1 => n2425, C2 => 
                           n1863, A => n1693, ZN => n1692);
   U1054 : AOI22_X1 port map( A1 => n1860, A2 => registers_17_31_port, B1 => 
                           n1859, B2 => registers_16_31_port, ZN => n1693);
   U1055 : OAI221_X1 port map( B1 => n1960, B2 => n2480, C1 => n1957, C2 => 
                           n2448, A => n715, ZN => n714);
   U1056 : AOI22_X1 port map( A1 => registers_17_8_port, A2 => n1954, B1 => 
                           registers_16_8_port, B2 => n1951, ZN => n715);
   U1057 : OAI221_X1 port map( B1 => n1960, B2 => n2479, C1 => n1957, C2 => 
                           n2447, A => n732, ZN => n731);
   U1058 : AOI22_X1 port map( A1 => registers_17_9_port, A2 => n1954, B1 => 
                           registers_16_9_port, B2 => n1951, ZN => n732);
   U1059 : OAI221_X1 port map( B1 => n1960, B2 => n2478, C1 => n1957, C2 => 
                           n2446, A => n749, ZN => n748);
   U1060 : AOI22_X1 port map( A1 => registers_17_10_port, A2 => n1954, B1 => 
                           registers_16_10_port, B2 => n1951, ZN => n749);
   U1061 : OAI221_X1 port map( B1 => n1960, B2 => n2477, C1 => n1957, C2 => 
                           n2445, A => n766, ZN => n765);
   U1062 : AOI22_X1 port map( A1 => registers_17_11_port, A2 => n1954, B1 => 
                           registers_16_11_port, B2 => n1951, ZN => n766);
   U1063 : OAI221_X1 port map( B1 => n1960, B2 => n2476, C1 => n1957, C2 => 
                           n2444, A => n783, ZN => n782);
   U1064 : AOI22_X1 port map( A1 => registers_17_12_port, A2 => n1954, B1 => 
                           registers_16_12_port, B2 => n1951, ZN => n783);
   U1065 : OAI221_X1 port map( B1 => n1960, B2 => n2475, C1 => n1957, C2 => 
                           n2443, A => n800, ZN => n799);
   U1066 : AOI22_X1 port map( A1 => registers_17_13_port, A2 => n1954, B1 => 
                           registers_16_13_port, B2 => n1951, ZN => n800);
   U1067 : OAI221_X1 port map( B1 => n1960, B2 => n2474, C1 => n1957, C2 => 
                           n2442, A => n817, ZN => n816);
   U1068 : AOI22_X1 port map( A1 => registers_17_14_port, A2 => n1954, B1 => 
                           registers_16_14_port, B2 => n1951, ZN => n817);
   U1069 : OAI221_X1 port map( B1 => n1960, B2 => n2473, C1 => n1957, C2 => 
                           n2441, A => n834, ZN => n833);
   U1070 : AOI22_X1 port map( A1 => registers_17_15_port, A2 => n1954, B1 => 
                           registers_16_15_port, B2 => n1951, ZN => n834);
   U1071 : OAI221_X1 port map( B1 => n1960, B2 => n2472, C1 => n1957, C2 => 
                           n2440, A => n851, ZN => n850);
   U1072 : AOI22_X1 port map( A1 => registers_17_16_port, A2 => n1954, B1 => 
                           registers_16_16_port, B2 => n1951, ZN => n851);
   U1073 : OAI221_X1 port map( B1 => n1960, B2 => n2471, C1 => n1957, C2 => 
                           n2439, A => n868, ZN => n867);
   U1074 : AOI22_X1 port map( A1 => registers_17_17_port, A2 => n1954, B1 => 
                           registers_16_17_port, B2 => n1951, ZN => n868);
   U1075 : OAI221_X1 port map( B1 => n1960, B2 => n2470, C1 => n1957, C2 => 
                           n2438, A => n885, ZN => n884);
   U1076 : AOI22_X1 port map( A1 => registers_17_18_port, A2 => n1954, B1 => 
                           registers_16_18_port, B2 => n1951, ZN => n885);
   U1077 : OAI221_X1 port map( B1 => n1960, B2 => n2469, C1 => n1957, C2 => 
                           n2437, A => n902, ZN => n901);
   U1078 : AOI22_X1 port map( A1 => registers_17_19_port, A2 => n1954, B1 => 
                           registers_16_19_port, B2 => n1951, ZN => n902);
   U1079 : OAI221_X1 port map( B1 => n1959, B2 => n2468, C1 => n1956, C2 => 
                           n2436, A => n919, ZN => n918);
   U1080 : AOI22_X1 port map( A1 => registers_17_20_port, A2 => n1953, B1 => 
                           registers_16_20_port, B2 => n1950, ZN => n919);
   U1081 : OAI221_X1 port map( B1 => n1959, B2 => n2467, C1 => n1956, C2 => 
                           n2435, A => n936, ZN => n935);
   U1082 : AOI22_X1 port map( A1 => registers_17_21_port, A2 => n1953, B1 => 
                           registers_16_21_port, B2 => n1950, ZN => n936);
   U1083 : OAI221_X1 port map( B1 => n1959, B2 => n2466, C1 => n1956, C2 => 
                           n2434, A => n953, ZN => n952);
   U1084 : AOI22_X1 port map( A1 => registers_17_22_port, A2 => n1953, B1 => 
                           registers_16_22_port, B2 => n1950, ZN => n953);
   U1085 : OAI221_X1 port map( B1 => n1959, B2 => n2465, C1 => n1956, C2 => 
                           n2433, A => n970, ZN => n969);
   U1086 : AOI22_X1 port map( A1 => registers_17_23_port, A2 => n1953, B1 => 
                           registers_16_23_port, B2 => n1950, ZN => n970);
   U1087 : OAI221_X1 port map( B1 => n1959, B2 => n2464, C1 => n1956, C2 => 
                           n2432, A => n987, ZN => n986);
   U1088 : AOI22_X1 port map( A1 => registers_17_24_port, A2 => n1953, B1 => 
                           registers_16_24_port, B2 => n1950, ZN => n987);
   U1089 : OAI221_X1 port map( B1 => n1959, B2 => n2463, C1 => n1956, C2 => 
                           n2431, A => n1004, ZN => n1003);
   U1090 : AOI22_X1 port map( A1 => registers_17_25_port, A2 => n1953, B1 => 
                           registers_16_25_port, B2 => n1950, ZN => n1004);
   U1091 : OAI221_X1 port map( B1 => n1959, B2 => n2462, C1 => n1956, C2 => 
                           n2430, A => n1021, ZN => n1020);
   U1092 : AOI22_X1 port map( A1 => registers_17_26_port, A2 => n1953, B1 => 
                           registers_16_26_port, B2 => n1950, ZN => n1021);
   U1093 : OAI221_X1 port map( B1 => n1959, B2 => n2461, C1 => n1956, C2 => 
                           n2429, A => n1038, ZN => n1037);
   U1094 : AOI22_X1 port map( A1 => registers_17_27_port, A2 => n1953, B1 => 
                           registers_16_27_port, B2 => n1950, ZN => n1038);
   U1095 : OAI221_X1 port map( B1 => n1959, B2 => n2460, C1 => n1956, C2 => 
                           n2428, A => n1055, ZN => n1054);
   U1096 : AOI22_X1 port map( A1 => registers_17_28_port, A2 => n1953, B1 => 
                           registers_16_28_port, B2 => n1950, ZN => n1055);
   U1097 : OAI221_X1 port map( B1 => n1959, B2 => n2459, C1 => n1956, C2 => 
                           n2427, A => n1072, ZN => n1071);
   U1098 : AOI22_X1 port map( A1 => registers_17_29_port, A2 => n1953, B1 => 
                           registers_16_29_port, B2 => n1950, ZN => n1072);
   U1099 : OAI221_X1 port map( B1 => n1959, B2 => n2458, C1 => n1956, C2 => 
                           n2426, A => n1089, ZN => n1088);
   U1100 : AOI22_X1 port map( A1 => registers_17_30_port, A2 => n1953, B1 => 
                           registers_16_30_port, B2 => n1950, ZN => n1089);
   U1101 : OAI221_X1 port map( B1 => n1959, B2 => n2457, C1 => n1956, C2 => 
                           n2425, A => n1106, ZN => n1105);
   U1102 : AOI22_X1 port map( A1 => registers_17_31_port, A2 => n1953, B1 => 
                           registers_16_31_port, B2 => n1950, ZN => n1106);
   U1103 : OAI221_X1 port map( B1 => n1904, B2 => n2200, C1 => n1901, C2 => 
                           n2264, A => n575, ZN => n569);
   U1104 : AOI22_X1 port map( A1 => registers_3_0_port, A2 => n1898, B1 => 
                           registers_6_0_port, B2 => n1895, ZN => n575);
   U1105 : OAI221_X1 port map( B1 => n1904, B2 => n2199, C1 => n1901, C2 => 
                           n2263, A => n602, ZN => n600);
   U1106 : AOI22_X1 port map( A1 => registers_3_1_port, A2 => n1898, B1 => 
                           registers_6_1_port, B2 => n1895, ZN => n602);
   U1107 : OAI221_X1 port map( B1 => n1904, B2 => n2198, C1 => n1901, C2 => 
                           n2262, A => n619, ZN => n617);
   U1108 : AOI22_X1 port map( A1 => registers_3_2_port, A2 => n1898, B1 => 
                           registers_6_2_port, B2 => n1895, ZN => n619);
   U1109 : OAI221_X1 port map( B1 => n1904, B2 => n2197, C1 => n1901, C2 => 
                           n2261, A => n636, ZN => n634);
   U1110 : AOI22_X1 port map( A1 => registers_3_3_port, A2 => n1898, B1 => 
                           registers_6_3_port, B2 => n1895, ZN => n636);
   U1111 : OAI221_X1 port map( B1 => n1904, B2 => n2196, C1 => n1901, C2 => 
                           n2260, A => n653, ZN => n651);
   U1112 : AOI22_X1 port map( A1 => registers_3_4_port, A2 => n1898, B1 => 
                           registers_6_4_port, B2 => n1895, ZN => n653);
   U1113 : OAI221_X1 port map( B1 => n1904, B2 => n2195, C1 => n1901, C2 => 
                           n2259, A => n670, ZN => n668);
   U1114 : AOI22_X1 port map( A1 => registers_3_5_port, A2 => n1898, B1 => 
                           registers_6_5_port, B2 => n1895, ZN => n670);
   U1115 : OAI221_X1 port map( B1 => n1904, B2 => n2194, C1 => n1901, C2 => 
                           n2258, A => n687, ZN => n685);
   U1116 : AOI22_X1 port map( A1 => registers_3_6_port, A2 => n1898, B1 => 
                           registers_6_6_port, B2 => n1895, ZN => n687);
   U1117 : OAI221_X1 port map( B1 => n1904, B2 => n2193, C1 => n1901, C2 => 
                           n2257, A => n704, ZN => n702);
   U1118 : AOI22_X1 port map( A1 => registers_3_7_port, A2 => n1898, B1 => 
                           registers_6_7_port, B2 => n1895, ZN => n704);
   U1119 : OAI221_X1 port map( B1 => n2200, B2 => n1811, C1 => n2264, C2 => 
                           n1808, A => n1162, ZN => n1156);
   U1120 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_0_port, B1 => 
                           n1800, B2 => registers_6_0_port, ZN => n1162);
   U1121 : OAI221_X1 port map( B1 => n2199, B2 => n1811, C1 => n2263, C2 => 
                           n1808, A => n1189, ZN => n1187);
   U1122 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_1_port, B1 => 
                           n1800, B2 => registers_6_1_port, ZN => n1189);
   U1123 : OAI221_X1 port map( B1 => n2198, B2 => n1811, C1 => n2262, C2 => 
                           n1808, A => n1206, ZN => n1204);
   U1124 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_2_port, B1 => 
                           n1800, B2 => registers_6_2_port, ZN => n1206);
   U1125 : OAI221_X1 port map( B1 => n2197, B2 => n1811, C1 => n2261, C2 => 
                           n1808, A => n1223, ZN => n1221);
   U1126 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_3_port, B1 => 
                           n1800, B2 => registers_6_3_port, ZN => n1223);
   U1127 : OAI221_X1 port map( B1 => n2196, B2 => n1811, C1 => n2260, C2 => 
                           n1808, A => n1240, ZN => n1238);
   U1128 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_4_port, B1 => 
                           n1800, B2 => registers_6_4_port, ZN => n1240);
   U1129 : OAI221_X1 port map( B1 => n2195, B2 => n1811, C1 => n2259, C2 => 
                           n1808, A => n1257, ZN => n1255);
   U1130 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_5_port, B1 => 
                           n1800, B2 => registers_6_5_port, ZN => n1257);
   U1131 : OAI221_X1 port map( B1 => n2194, B2 => n1811, C1 => n2258, C2 => 
                           n1808, A => n1274, ZN => n1272);
   U1132 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_6_port, B1 => 
                           n1800, B2 => registers_6_6_port, ZN => n1274);
   U1133 : OAI221_X1 port map( B1 => n2193, B2 => n1811, C1 => n2257, C2 => 
                           n1808, A => n1291, ZN => n1289);
   U1134 : AOI22_X1 port map( A1 => n1805, A2 => registers_3_7_port, B1 => 
                           n1800, B2 => registers_6_7_port, ZN => n1291);
   U1135 : OAI221_X1 port map( B1 => n2192, B2 => n1810, C1 => n2256, C2 => 
                           n1807, A => n1308, ZN => n1306);
   U1136 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_8_port, B1 => 
                           n1800, B2 => registers_6_8_port, ZN => n1308);
   U1137 : OAI221_X1 port map( B1 => n2191, B2 => n1810, C1 => n2255, C2 => 
                           n1807, A => n1325, ZN => n1323);
   U1138 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_9_port, B1 => 
                           n1800, B2 => registers_6_9_port, ZN => n1325);
   U1139 : OAI221_X1 port map( B1 => n2190, B2 => n1810, C1 => n2254, C2 => 
                           n1807, A => n1342, ZN => n1340);
   U1140 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_10_port, B1 => 
                           n1800, B2 => registers_6_10_port, ZN => n1342);
   U1141 : OAI221_X1 port map( B1 => n2189, B2 => n1810, C1 => n2253, C2 => 
                           n1807, A => n1359, ZN => n1357);
   U1142 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_11_port, B1 => 
                           n1800, B2 => registers_6_11_port, ZN => n1359);
   U1143 : OAI221_X1 port map( B1 => n2188, B2 => n1810, C1 => n2252, C2 => 
                           n1807, A => n1376, ZN => n1374);
   U1144 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_12_port, B1 => 
                           n1801, B2 => registers_6_12_port, ZN => n1376);
   U1145 : OAI221_X1 port map( B1 => n2187, B2 => n1810, C1 => n2251, C2 => 
                           n1807, A => n1393, ZN => n1391);
   U1146 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_13_port, B1 => 
                           n1801, B2 => registers_6_13_port, ZN => n1393);
   U1147 : OAI221_X1 port map( B1 => n2186, B2 => n1810, C1 => n2250, C2 => 
                           n1807, A => n1410, ZN => n1408);
   U1148 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_14_port, B1 => 
                           n1801, B2 => registers_6_14_port, ZN => n1410);
   U1149 : OAI221_X1 port map( B1 => n2185, B2 => n1810, C1 => n2249, C2 => 
                           n1807, A => n1427, ZN => n1425);
   U1150 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_15_port, B1 => 
                           n1801, B2 => registers_6_15_port, ZN => n1427);
   U1151 : OAI221_X1 port map( B1 => n2184, B2 => n1810, C1 => n2248, C2 => 
                           n1807, A => n1444, ZN => n1442);
   U1152 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_16_port, B1 => 
                           n1801, B2 => registers_6_16_port, ZN => n1444);
   U1153 : OAI221_X1 port map( B1 => n2183, B2 => n1810, C1 => n2247, C2 => 
                           n1807, A => n1461, ZN => n1459);
   U1154 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_17_port, B1 => 
                           n1801, B2 => registers_6_17_port, ZN => n1461);
   U1155 : OAI221_X1 port map( B1 => n2182, B2 => n1810, C1 => n2246, C2 => 
                           n1807, A => n1478, ZN => n1476);
   U1156 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_18_port, B1 => 
                           n1801, B2 => registers_6_18_port, ZN => n1478);
   U1157 : OAI221_X1 port map( B1 => n2181, B2 => n1810, C1 => n2245, C2 => 
                           n1807, A => n1495, ZN => n1493);
   U1158 : AOI22_X1 port map( A1 => n1804, A2 => registers_3_19_port, B1 => 
                           n1801, B2 => registers_6_19_port, ZN => n1495);
   U1159 : OAI221_X1 port map( B1 => n2180, B2 => n1809, C1 => n2244, C2 => 
                           n1806, A => n1512, ZN => n1510);
   U1160 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_20_port, B1 => 
                           n1801, B2 => registers_6_20_port, ZN => n1512);
   U1161 : OAI221_X1 port map( B1 => n2179, B2 => n1809, C1 => n2243, C2 => 
                           n1806, A => n1529, ZN => n1527);
   U1162 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_21_port, B1 => 
                           n1801, B2 => registers_6_21_port, ZN => n1529);
   U1163 : OAI221_X1 port map( B1 => n2178, B2 => n1809, C1 => n2242, C2 => 
                           n1806, A => n1546, ZN => n1544);
   U1164 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_22_port, B1 => 
                           n1801, B2 => registers_6_22_port, ZN => n1546);
   U1165 : OAI221_X1 port map( B1 => n2177, B2 => n1809, C1 => n2241, C2 => 
                           n1806, A => n1563, ZN => n1561);
   U1166 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_23_port, B1 => 
                           n1801, B2 => registers_6_23_port, ZN => n1563);
   U1167 : OAI221_X1 port map( B1 => n2176, B2 => n1809, C1 => n2240, C2 => 
                           n1806, A => n1580, ZN => n1578);
   U1168 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_24_port, B1 => 
                           n1802, B2 => registers_6_24_port, ZN => n1580);
   U1169 : OAI221_X1 port map( B1 => n2175, B2 => n1809, C1 => n2239, C2 => 
                           n1806, A => n1597, ZN => n1595);
   U1170 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_25_port, B1 => 
                           n1802, B2 => registers_6_25_port, ZN => n1597);
   U1171 : OAI221_X1 port map( B1 => n2174, B2 => n1809, C1 => n2238, C2 => 
                           n1806, A => n1614, ZN => n1612);
   U1172 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_26_port, B1 => 
                           n1802, B2 => registers_6_26_port, ZN => n1614);
   U1173 : OAI221_X1 port map( B1 => n2173, B2 => n1809, C1 => n2237, C2 => 
                           n1806, A => n1631, ZN => n1629);
   U1174 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_27_port, B1 => 
                           n1802, B2 => registers_6_27_port, ZN => n1631);
   U1175 : OAI221_X1 port map( B1 => n2172, B2 => n1809, C1 => n2236, C2 => 
                           n1806, A => n1648, ZN => n1646);
   U1176 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_28_port, B1 => 
                           n1802, B2 => registers_6_28_port, ZN => n1648);
   U1177 : OAI221_X1 port map( B1 => n2171, B2 => n1809, C1 => n2235, C2 => 
                           n1806, A => n1665, ZN => n1663);
   U1178 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_29_port, B1 => 
                           n1802, B2 => registers_6_29_port, ZN => n1665);
   U1179 : OAI221_X1 port map( B1 => n2170, B2 => n1809, C1 => n2234, C2 => 
                           n1806, A => n1682, ZN => n1680);
   U1180 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_30_port, B1 => 
                           n1802, B2 => registers_6_30_port, ZN => n1682);
   U1181 : OAI221_X1 port map( B1 => n2169, B2 => n1809, C1 => n2233, C2 => 
                           n1806, A => n1709, ZN => n1705);
   U1182 : AOI22_X1 port map( A1 => n1803, A2 => registers_3_31_port, B1 => 
                           n1802, B2 => registers_6_31_port, ZN => n1709);
   U1183 : OAI221_X1 port map( B1 => n1903, B2 => n2192, C1 => n1900, C2 => 
                           n2256, A => n721, ZN => n719);
   U1184 : AOI22_X1 port map( A1 => registers_3_8_port, A2 => n1897, B1 => 
                           registers_6_8_port, B2 => n1894, ZN => n721);
   U1185 : OAI221_X1 port map( B1 => n1903, B2 => n2191, C1 => n1900, C2 => 
                           n2255, A => n738, ZN => n736);
   U1186 : AOI22_X1 port map( A1 => registers_3_9_port, A2 => n1897, B1 => 
                           registers_6_9_port, B2 => n1894, ZN => n738);
   U1187 : OAI221_X1 port map( B1 => n1903, B2 => n2190, C1 => n1900, C2 => 
                           n2254, A => n755, ZN => n753);
   U1188 : AOI22_X1 port map( A1 => registers_3_10_port, A2 => n1897, B1 => 
                           registers_6_10_port, B2 => n1894, ZN => n755);
   U1189 : OAI221_X1 port map( B1 => n1903, B2 => n2189, C1 => n1900, C2 => 
                           n2253, A => n772, ZN => n770);
   U1190 : AOI22_X1 port map( A1 => registers_3_11_port, A2 => n1897, B1 => 
                           registers_6_11_port, B2 => n1894, ZN => n772);
   U1191 : OAI221_X1 port map( B1 => n1903, B2 => n2188, C1 => n1900, C2 => 
                           n2252, A => n789, ZN => n787);
   U1192 : AOI22_X1 port map( A1 => registers_3_12_port, A2 => n1897, B1 => 
                           registers_6_12_port, B2 => n1894, ZN => n789);
   U1193 : OAI221_X1 port map( B1 => n1903, B2 => n2187, C1 => n1900, C2 => 
                           n2251, A => n806, ZN => n804);
   U1194 : AOI22_X1 port map( A1 => registers_3_13_port, A2 => n1897, B1 => 
                           registers_6_13_port, B2 => n1894, ZN => n806);
   U1195 : OAI221_X1 port map( B1 => n1903, B2 => n2186, C1 => n1900, C2 => 
                           n2250, A => n823, ZN => n821);
   U1196 : AOI22_X1 port map( A1 => registers_3_14_port, A2 => n1897, B1 => 
                           registers_6_14_port, B2 => n1894, ZN => n823);
   U1197 : OAI221_X1 port map( B1 => n1903, B2 => n2185, C1 => n1900, C2 => 
                           n2249, A => n840, ZN => n838);
   U1198 : AOI22_X1 port map( A1 => registers_3_15_port, A2 => n1897, B1 => 
                           registers_6_15_port, B2 => n1894, ZN => n840);
   U1199 : OAI221_X1 port map( B1 => n1903, B2 => n2184, C1 => n1900, C2 => 
                           n2248, A => n857, ZN => n855);
   U1200 : AOI22_X1 port map( A1 => registers_3_16_port, A2 => n1897, B1 => 
                           registers_6_16_port, B2 => n1894, ZN => n857);
   U1201 : OAI221_X1 port map( B1 => n1903, B2 => n2183, C1 => n1900, C2 => 
                           n2247, A => n874, ZN => n872);
   U1202 : AOI22_X1 port map( A1 => registers_3_17_port, A2 => n1897, B1 => 
                           registers_6_17_port, B2 => n1894, ZN => n874);
   U1203 : OAI221_X1 port map( B1 => n1903, B2 => n2182, C1 => n1900, C2 => 
                           n2246, A => n891, ZN => n889);
   U1204 : AOI22_X1 port map( A1 => registers_3_18_port, A2 => n1897, B1 => 
                           registers_6_18_port, B2 => n1894, ZN => n891);
   U1205 : OAI221_X1 port map( B1 => n1903, B2 => n2181, C1 => n1900, C2 => 
                           n2245, A => n908, ZN => n906);
   U1206 : AOI22_X1 port map( A1 => registers_3_19_port, A2 => n1897, B1 => 
                           registers_6_19_port, B2 => n1894, ZN => n908);
   U1207 : OAI221_X1 port map( B1 => n1902, B2 => n2180, C1 => n1899, C2 => 
                           n2244, A => n925, ZN => n923);
   U1208 : AOI22_X1 port map( A1 => registers_3_20_port, A2 => n1896, B1 => 
                           registers_6_20_port, B2 => n1893, ZN => n925);
   U1209 : OAI221_X1 port map( B1 => n1902, B2 => n2179, C1 => n1899, C2 => 
                           n2243, A => n942, ZN => n940);
   U1210 : AOI22_X1 port map( A1 => registers_3_21_port, A2 => n1896, B1 => 
                           registers_6_21_port, B2 => n1893, ZN => n942);
   U1211 : OAI221_X1 port map( B1 => n1902, B2 => n2178, C1 => n1899, C2 => 
                           n2242, A => n959, ZN => n957);
   U1212 : AOI22_X1 port map( A1 => registers_3_22_port, A2 => n1896, B1 => 
                           registers_6_22_port, B2 => n1893, ZN => n959);
   U1213 : OAI221_X1 port map( B1 => n1902, B2 => n2177, C1 => n1899, C2 => 
                           n2241, A => n976, ZN => n974);
   U1214 : AOI22_X1 port map( A1 => registers_3_23_port, A2 => n1896, B1 => 
                           registers_6_23_port, B2 => n1893, ZN => n976);
   U1215 : OAI221_X1 port map( B1 => n1902, B2 => n2176, C1 => n1899, C2 => 
                           n2240, A => n993, ZN => n991);
   U1216 : AOI22_X1 port map( A1 => registers_3_24_port, A2 => n1896, B1 => 
                           registers_6_24_port, B2 => n1893, ZN => n993);
   U1217 : OAI221_X1 port map( B1 => n1902, B2 => n2175, C1 => n1899, C2 => 
                           n2239, A => n1010, ZN => n1008);
   U1218 : AOI22_X1 port map( A1 => registers_3_25_port, A2 => n1896, B1 => 
                           registers_6_25_port, B2 => n1893, ZN => n1010);
   U1219 : OAI221_X1 port map( B1 => n1902, B2 => n2174, C1 => n1899, C2 => 
                           n2238, A => n1027, ZN => n1025);
   U1220 : AOI22_X1 port map( A1 => registers_3_26_port, A2 => n1896, B1 => 
                           registers_6_26_port, B2 => n1893, ZN => n1027);
   U1221 : OAI221_X1 port map( B1 => n1902, B2 => n2173, C1 => n1899, C2 => 
                           n2237, A => n1044, ZN => n1042);
   U1222 : AOI22_X1 port map( A1 => registers_3_27_port, A2 => n1896, B1 => 
                           registers_6_27_port, B2 => n1893, ZN => n1044);
   U1223 : OAI221_X1 port map( B1 => n1902, B2 => n2172, C1 => n1899, C2 => 
                           n2236, A => n1061, ZN => n1059);
   U1224 : AOI22_X1 port map( A1 => registers_3_28_port, A2 => n1896, B1 => 
                           registers_6_28_port, B2 => n1893, ZN => n1061);
   U1225 : OAI221_X1 port map( B1 => n1902, B2 => n2171, C1 => n1899, C2 => 
                           n2235, A => n1078, ZN => n1076);
   U1226 : AOI22_X1 port map( A1 => registers_3_29_port, A2 => n1896, B1 => 
                           registers_6_29_port, B2 => n1893, ZN => n1078);
   U1227 : OAI221_X1 port map( B1 => n1902, B2 => n2170, C1 => n1899, C2 => 
                           n2234, A => n1095, ZN => n1093);
   U1228 : AOI22_X1 port map( A1 => registers_3_30_port, A2 => n1896, B1 => 
                           registers_6_30_port, B2 => n1893, ZN => n1095);
   U1229 : OAI221_X1 port map( B1 => n1902, B2 => n2169, C1 => n1899, C2 => 
                           n2233, A => n1122, ZN => n1118);
   U1230 : AOI22_X1 port map( A1 => registers_3_31_port, A2 => n1896, B1 => 
                           registers_6_31_port, B2 => n1893, ZN => n1122);
   U1231 : AOI22_X1 port map( A1 => registers_23_0_port, A2 => n1943, B1 => 
                           registers_22_0_port, B2 => n1940, ZN => n555);
   U1232 : AOI22_X1 port map( A1 => registers_25_0_port, A2 => n1931, B1 => 
                           registers_24_0_port, B2 => n1928, ZN => n560);
   U1233 : AOI22_X1 port map( A1 => registers_31_0_port, A2 => n1919, B1 => 
                           registers_30_0_port, B2 => n1916, ZN => n565);
   U1234 : AOI22_X1 port map( A1 => registers_23_1_port, A2 => n1943, B1 => 
                           registers_22_1_port, B2 => n1940, ZN => n597);
   U1235 : AOI22_X1 port map( A1 => registers_25_1_port, A2 => n1931, B1 => 
                           registers_24_1_port, B2 => n1928, ZN => n598);
   U1236 : AOI22_X1 port map( A1 => registers_31_1_port, A2 => n1919, B1 => 
                           registers_30_1_port, B2 => n1916, ZN => n599);
   U1237 : AOI22_X1 port map( A1 => registers_23_2_port, A2 => n1943, B1 => 
                           registers_22_2_port, B2 => n1940, ZN => n614);
   U1238 : AOI22_X1 port map( A1 => registers_25_2_port, A2 => n1931, B1 => 
                           registers_24_2_port, B2 => n1928, ZN => n615);
   U1239 : AOI22_X1 port map( A1 => registers_31_2_port, A2 => n1919, B1 => 
                           registers_30_2_port, B2 => n1916, ZN => n616);
   U1240 : AOI22_X1 port map( A1 => registers_23_3_port, A2 => n1943, B1 => 
                           registers_22_3_port, B2 => n1940, ZN => n631);
   U1241 : AOI22_X1 port map( A1 => registers_25_3_port, A2 => n1931, B1 => 
                           registers_24_3_port, B2 => n1928, ZN => n632);
   U1242 : AOI22_X1 port map( A1 => registers_31_3_port, A2 => n1919, B1 => 
                           registers_30_3_port, B2 => n1916, ZN => n633);
   U1243 : AOI22_X1 port map( A1 => registers_23_4_port, A2 => n1943, B1 => 
                           registers_22_4_port, B2 => n1940, ZN => n648);
   U1244 : AOI22_X1 port map( A1 => registers_25_4_port, A2 => n1931, B1 => 
                           registers_24_4_port, B2 => n1928, ZN => n649);
   U1245 : AOI22_X1 port map( A1 => registers_31_4_port, A2 => n1919, B1 => 
                           registers_30_4_port, B2 => n1916, ZN => n650);
   U1246 : AOI22_X1 port map( A1 => registers_23_5_port, A2 => n1943, B1 => 
                           registers_22_5_port, B2 => n1940, ZN => n665);
   U1247 : AOI22_X1 port map( A1 => registers_25_5_port, A2 => n1931, B1 => 
                           registers_24_5_port, B2 => n1928, ZN => n666);
   U1248 : AOI22_X1 port map( A1 => registers_31_5_port, A2 => n1919, B1 => 
                           registers_30_5_port, B2 => n1916, ZN => n667);
   U1249 : AOI22_X1 port map( A1 => registers_23_6_port, A2 => n1943, B1 => 
                           registers_22_6_port, B2 => n1940, ZN => n682);
   U1250 : AOI22_X1 port map( A1 => registers_25_6_port, A2 => n1931, B1 => 
                           registers_24_6_port, B2 => n1928, ZN => n683);
   U1251 : AOI22_X1 port map( A1 => registers_31_6_port, A2 => n1919, B1 => 
                           registers_30_6_port, B2 => n1916, ZN => n684);
   U1252 : AOI22_X1 port map( A1 => registers_23_7_port, A2 => n1943, B1 => 
                           registers_22_7_port, B2 => n1940, ZN => n699);
   U1253 : AOI22_X1 port map( A1 => registers_25_7_port, A2 => n1931, B1 => 
                           registers_24_7_port, B2 => n1928, ZN => n700);
   U1254 : AOI22_X1 port map( A1 => registers_31_7_port, A2 => n1919, B1 => 
                           registers_30_7_port, B2 => n1916, ZN => n701);
   U1255 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_0_port, B1 => 
                           n1845, B2 => registers_22_0_port, ZN => n1142);
   U1256 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_0_port, B1 => 
                           n1833, B2 => registers_24_0_port, ZN => n1147);
   U1257 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_0_port, B1 => 
                           n1821, B2 => registers_30_0_port, ZN => n1152);
   U1258 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_1_port, B1 => 
                           n1845, B2 => registers_22_1_port, ZN => n1184);
   U1259 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_1_port, B1 => 
                           n1833, B2 => registers_24_1_port, ZN => n1185);
   U1260 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_1_port, B1 => 
                           n1821, B2 => registers_30_1_port, ZN => n1186);
   U1261 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_2_port, B1 => 
                           n1845, B2 => registers_22_2_port, ZN => n1201);
   U1262 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_2_port, B1 => 
                           n1833, B2 => registers_24_2_port, ZN => n1202);
   U1263 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_2_port, B1 => 
                           n1821, B2 => registers_30_2_port, ZN => n1203);
   U1264 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_3_port, B1 => 
                           n1845, B2 => registers_22_3_port, ZN => n1218);
   U1265 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_3_port, B1 => 
                           n1833, B2 => registers_24_3_port, ZN => n1219);
   U1266 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_3_port, B1 => 
                           n1821, B2 => registers_30_3_port, ZN => n1220);
   U1267 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_4_port, B1 => 
                           n1845, B2 => registers_22_4_port, ZN => n1235);
   U1268 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_4_port, B1 => 
                           n1833, B2 => registers_24_4_port, ZN => n1236);
   U1269 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_4_port, B1 => 
                           n1821, B2 => registers_30_4_port, ZN => n1237);
   U1270 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_5_port, B1 => 
                           n1845, B2 => registers_22_5_port, ZN => n1252);
   U1271 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_5_port, B1 => 
                           n1833, B2 => registers_24_5_port, ZN => n1253);
   U1272 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_5_port, B1 => 
                           n1821, B2 => registers_30_5_port, ZN => n1254);
   U1273 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_6_port, B1 => 
                           n1845, B2 => registers_22_6_port, ZN => n1269);
   U1274 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_6_port, B1 => 
                           n1833, B2 => registers_24_6_port, ZN => n1270);
   U1275 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_6_port, B1 => 
                           n1821, B2 => registers_30_6_port, ZN => n1271);
   U1276 : AOI22_X1 port map( A1 => n1850, A2 => registers_23_7_port, B1 => 
                           n1845, B2 => registers_22_7_port, ZN => n1286);
   U1277 : AOI22_X1 port map( A1 => n1838, A2 => registers_25_7_port, B1 => 
                           n1833, B2 => registers_24_7_port, ZN => n1287);
   U1278 : AOI22_X1 port map( A1 => n1826, A2 => registers_31_7_port, B1 => 
                           n1821, B2 => registers_30_7_port, ZN => n1288);
   U1279 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_8_port, B1 => 
                           n1845, B2 => registers_22_8_port, ZN => n1303);
   U1280 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_8_port, B1 => 
                           n1833, B2 => registers_24_8_port, ZN => n1304);
   U1281 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_8_port, B1 => 
                           n1821, B2 => registers_30_8_port, ZN => n1305);
   U1282 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_9_port, B1 => 
                           n1845, B2 => registers_22_9_port, ZN => n1320);
   U1283 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_9_port, B1 => 
                           n1833, B2 => registers_24_9_port, ZN => n1321);
   U1284 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_9_port, B1 => 
                           n1821, B2 => registers_30_9_port, ZN => n1322);
   U1285 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_10_port, B1 => 
                           n1845, B2 => registers_22_10_port, ZN => n1337);
   U1286 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_10_port, B1 => 
                           n1833, B2 => registers_24_10_port, ZN => n1338);
   U1287 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_10_port, B1 => 
                           n1821, B2 => registers_30_10_port, ZN => n1339);
   U1288 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_11_port, B1 => 
                           n1845, B2 => registers_22_11_port, ZN => n1354);
   U1289 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_11_port, B1 => 
                           n1833, B2 => registers_24_11_port, ZN => n1355);
   U1290 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_11_port, B1 => 
                           n1821, B2 => registers_30_11_port, ZN => n1356);
   U1291 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_12_port, B1 => 
                           n1846, B2 => registers_22_12_port, ZN => n1371);
   U1292 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_12_port, B1 => 
                           n1834, B2 => registers_24_12_port, ZN => n1372);
   U1293 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_12_port, B1 => 
                           n1822, B2 => registers_30_12_port, ZN => n1373);
   U1294 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_13_port, B1 => 
                           n1846, B2 => registers_22_13_port, ZN => n1388);
   U1295 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_13_port, B1 => 
                           n1834, B2 => registers_24_13_port, ZN => n1389);
   U1296 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_13_port, B1 => 
                           n1822, B2 => registers_30_13_port, ZN => n1390);
   U1297 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_14_port, B1 => 
                           n1846, B2 => registers_22_14_port, ZN => n1405);
   U1298 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_14_port, B1 => 
                           n1834, B2 => registers_24_14_port, ZN => n1406);
   U1299 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_14_port, B1 => 
                           n1822, B2 => registers_30_14_port, ZN => n1407);
   U1300 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_15_port, B1 => 
                           n1846, B2 => registers_22_15_port, ZN => n1422);
   U1301 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_15_port, B1 => 
                           n1834, B2 => registers_24_15_port, ZN => n1423);
   U1302 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_15_port, B1 => 
                           n1822, B2 => registers_30_15_port, ZN => n1424);
   U1303 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_16_port, B1 => 
                           n1846, B2 => registers_22_16_port, ZN => n1439);
   U1304 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_16_port, B1 => 
                           n1834, B2 => registers_24_16_port, ZN => n1440);
   U1305 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_16_port, B1 => 
                           n1822, B2 => registers_30_16_port, ZN => n1441);
   U1306 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_17_port, B1 => 
                           n1846, B2 => registers_22_17_port, ZN => n1456);
   U1307 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_17_port, B1 => 
                           n1834, B2 => registers_24_17_port, ZN => n1457);
   U1308 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_17_port, B1 => 
                           n1822, B2 => registers_30_17_port, ZN => n1458);
   U1309 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_18_port, B1 => 
                           n1846, B2 => registers_22_18_port, ZN => n1473);
   U1310 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_18_port, B1 => 
                           n1834, B2 => registers_24_18_port, ZN => n1474);
   U1311 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_18_port, B1 => 
                           n1822, B2 => registers_30_18_port, ZN => n1475);
   U1312 : AOI22_X1 port map( A1 => n1849, A2 => registers_23_19_port, B1 => 
                           n1846, B2 => registers_22_19_port, ZN => n1490);
   U1313 : AOI22_X1 port map( A1 => n1837, A2 => registers_25_19_port, B1 => 
                           n1834, B2 => registers_24_19_port, ZN => n1491);
   U1314 : AOI22_X1 port map( A1 => n1825, A2 => registers_31_19_port, B1 => 
                           n1822, B2 => registers_30_19_port, ZN => n1492);
   U1315 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_20_port, B1 => 
                           n1846, B2 => registers_22_20_port, ZN => n1507);
   U1316 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_20_port, B1 => 
                           n1834, B2 => registers_24_20_port, ZN => n1508);
   U1317 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_20_port, B1 => 
                           n1822, B2 => registers_30_20_port, ZN => n1509);
   U1318 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_21_port, B1 => 
                           n1846, B2 => registers_22_21_port, ZN => n1524);
   U1319 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_21_port, B1 => 
                           n1834, B2 => registers_24_21_port, ZN => n1525);
   U1320 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_21_port, B1 => 
                           n1822, B2 => registers_30_21_port, ZN => n1526);
   U1321 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_22_port, B1 => 
                           n1846, B2 => registers_22_22_port, ZN => n1541);
   U1322 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_22_port, B1 => 
                           n1834, B2 => registers_24_22_port, ZN => n1542);
   U1323 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_22_port, B1 => 
                           n1822, B2 => registers_30_22_port, ZN => n1543);
   U1324 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_23_port, B1 => 
                           n1846, B2 => registers_22_23_port, ZN => n1558);
   U1325 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_23_port, B1 => 
                           n1834, B2 => registers_24_23_port, ZN => n1559);
   U1326 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_23_port, B1 => 
                           n1822, B2 => registers_30_23_port, ZN => n1560);
   U1327 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_24_port, B1 => 
                           n1847, B2 => registers_22_24_port, ZN => n1575);
   U1328 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_24_port, B1 => 
                           n1835, B2 => registers_24_24_port, ZN => n1576);
   U1329 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_24_port, B1 => 
                           n1823, B2 => registers_30_24_port, ZN => n1577);
   U1330 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_25_port, B1 => 
                           n1847, B2 => registers_22_25_port, ZN => n1592);
   U1331 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_25_port, B1 => 
                           n1835, B2 => registers_24_25_port, ZN => n1593);
   U1332 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_25_port, B1 => 
                           n1823, B2 => registers_30_25_port, ZN => n1594);
   U1333 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_26_port, B1 => 
                           n1847, B2 => registers_22_26_port, ZN => n1609);
   U1334 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_26_port, B1 => 
                           n1835, B2 => registers_24_26_port, ZN => n1610);
   U1335 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_26_port, B1 => 
                           n1823, B2 => registers_30_26_port, ZN => n1611);
   U1336 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_27_port, B1 => 
                           n1847, B2 => registers_22_27_port, ZN => n1626);
   U1337 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_27_port, B1 => 
                           n1835, B2 => registers_24_27_port, ZN => n1627);
   U1338 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_27_port, B1 => 
                           n1823, B2 => registers_30_27_port, ZN => n1628);
   U1339 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_28_port, B1 => 
                           n1847, B2 => registers_22_28_port, ZN => n1643);
   U1340 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_28_port, B1 => 
                           n1835, B2 => registers_24_28_port, ZN => n1644);
   U1341 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_28_port, B1 => 
                           n1823, B2 => registers_30_28_port, ZN => n1645);
   U1342 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_29_port, B1 => 
                           n1847, B2 => registers_22_29_port, ZN => n1660);
   U1343 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_29_port, B1 => 
                           n1835, B2 => registers_24_29_port, ZN => n1661);
   U1344 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_29_port, B1 => 
                           n1823, B2 => registers_30_29_port, ZN => n1662);
   U1345 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_30_port, B1 => 
                           n1847, B2 => registers_22_30_port, ZN => n1677);
   U1346 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_30_port, B1 => 
                           n1835, B2 => registers_24_30_port, ZN => n1678);
   U1347 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_30_port, B1 => 
                           n1823, B2 => registers_30_30_port, ZN => n1679);
   U1348 : AOI22_X1 port map( A1 => n1848, A2 => registers_23_31_port, B1 => 
                           n1847, B2 => registers_22_31_port, ZN => n1698);
   U1349 : AOI22_X1 port map( A1 => n1836, A2 => registers_25_31_port, B1 => 
                           n1835, B2 => registers_24_31_port, ZN => n1701);
   U1350 : AOI22_X1 port map( A1 => n1824, A2 => registers_31_31_port, B1 => 
                           n1823, B2 => registers_30_31_port, ZN => n1704);
   U1351 : AOI22_X1 port map( A1 => registers_23_8_port, A2 => n1942, B1 => 
                           registers_22_8_port, B2 => n1939, ZN => n716);
   U1352 : AOI22_X1 port map( A1 => registers_25_8_port, A2 => n1930, B1 => 
                           registers_24_8_port, B2 => n1927, ZN => n717);
   U1353 : AOI22_X1 port map( A1 => registers_31_8_port, A2 => n1918, B1 => 
                           registers_30_8_port, B2 => n1915, ZN => n718);
   U1354 : AOI22_X1 port map( A1 => registers_23_9_port, A2 => n1942, B1 => 
                           registers_22_9_port, B2 => n1939, ZN => n733);
   U1355 : AOI22_X1 port map( A1 => registers_25_9_port, A2 => n1930, B1 => 
                           registers_24_9_port, B2 => n1927, ZN => n734);
   U1356 : AOI22_X1 port map( A1 => registers_31_9_port, A2 => n1918, B1 => 
                           registers_30_9_port, B2 => n1915, ZN => n735);
   U1357 : AOI22_X1 port map( A1 => registers_23_10_port, A2 => n1942, B1 => 
                           registers_22_10_port, B2 => n1939, ZN => n750);
   U1358 : AOI22_X1 port map( A1 => registers_25_10_port, A2 => n1930, B1 => 
                           registers_24_10_port, B2 => n1927, ZN => n751);
   U1359 : AOI22_X1 port map( A1 => registers_31_10_port, A2 => n1918, B1 => 
                           registers_30_10_port, B2 => n1915, ZN => n752);
   U1360 : AOI22_X1 port map( A1 => registers_23_11_port, A2 => n1942, B1 => 
                           registers_22_11_port, B2 => n1939, ZN => n767);
   U1361 : AOI22_X1 port map( A1 => registers_25_11_port, A2 => n1930, B1 => 
                           registers_24_11_port, B2 => n1927, ZN => n768);
   U1362 : AOI22_X1 port map( A1 => registers_31_11_port, A2 => n1918, B1 => 
                           registers_30_11_port, B2 => n1915, ZN => n769);
   U1363 : AOI22_X1 port map( A1 => registers_23_12_port, A2 => n1942, B1 => 
                           registers_22_12_port, B2 => n1939, ZN => n784);
   U1364 : AOI22_X1 port map( A1 => registers_25_12_port, A2 => n1930, B1 => 
                           registers_24_12_port, B2 => n1927, ZN => n785);
   U1365 : AOI22_X1 port map( A1 => registers_31_12_port, A2 => n1918, B1 => 
                           registers_30_12_port, B2 => n1915, ZN => n786);
   U1366 : AOI22_X1 port map( A1 => registers_23_13_port, A2 => n1942, B1 => 
                           registers_22_13_port, B2 => n1939, ZN => n801);
   U1367 : AOI22_X1 port map( A1 => registers_25_13_port, A2 => n1930, B1 => 
                           registers_24_13_port, B2 => n1927, ZN => n802);
   U1368 : AOI22_X1 port map( A1 => registers_31_13_port, A2 => n1918, B1 => 
                           registers_30_13_port, B2 => n1915, ZN => n803);
   U1369 : AOI22_X1 port map( A1 => registers_23_14_port, A2 => n1942, B1 => 
                           registers_22_14_port, B2 => n1939, ZN => n818);
   U1370 : AOI22_X1 port map( A1 => registers_25_14_port, A2 => n1930, B1 => 
                           registers_24_14_port, B2 => n1927, ZN => n819);
   U1371 : AOI22_X1 port map( A1 => registers_31_14_port, A2 => n1918, B1 => 
                           registers_30_14_port, B2 => n1915, ZN => n820);
   U1372 : AOI22_X1 port map( A1 => registers_23_15_port, A2 => n1942, B1 => 
                           registers_22_15_port, B2 => n1939, ZN => n835);
   U1373 : AOI22_X1 port map( A1 => registers_25_15_port, A2 => n1930, B1 => 
                           registers_24_15_port, B2 => n1927, ZN => n836);
   U1374 : AOI22_X1 port map( A1 => registers_31_15_port, A2 => n1918, B1 => 
                           registers_30_15_port, B2 => n1915, ZN => n837);
   U1375 : AOI22_X1 port map( A1 => registers_23_16_port, A2 => n1942, B1 => 
                           registers_22_16_port, B2 => n1939, ZN => n852);
   U1376 : AOI22_X1 port map( A1 => registers_25_16_port, A2 => n1930, B1 => 
                           registers_24_16_port, B2 => n1927, ZN => n853);
   U1377 : AOI22_X1 port map( A1 => registers_31_16_port, A2 => n1918, B1 => 
                           registers_30_16_port, B2 => n1915, ZN => n854);
   U1378 : AOI22_X1 port map( A1 => registers_23_17_port, A2 => n1942, B1 => 
                           registers_22_17_port, B2 => n1939, ZN => n869);
   U1379 : AOI22_X1 port map( A1 => registers_25_17_port, A2 => n1930, B1 => 
                           registers_24_17_port, B2 => n1927, ZN => n870);
   U1380 : AOI22_X1 port map( A1 => registers_31_17_port, A2 => n1918, B1 => 
                           registers_30_17_port, B2 => n1915, ZN => n871);
   U1381 : AOI22_X1 port map( A1 => registers_23_18_port, A2 => n1942, B1 => 
                           registers_22_18_port, B2 => n1939, ZN => n886);
   U1382 : AOI22_X1 port map( A1 => registers_25_18_port, A2 => n1930, B1 => 
                           registers_24_18_port, B2 => n1927, ZN => n887);
   U1383 : AOI22_X1 port map( A1 => registers_31_18_port, A2 => n1918, B1 => 
                           registers_30_18_port, B2 => n1915, ZN => n888);
   U1384 : AOI22_X1 port map( A1 => registers_23_19_port, A2 => n1942, B1 => 
                           registers_22_19_port, B2 => n1939, ZN => n903);
   U1385 : AOI22_X1 port map( A1 => registers_25_19_port, A2 => n1930, B1 => 
                           registers_24_19_port, B2 => n1927, ZN => n904);
   U1386 : AOI22_X1 port map( A1 => registers_31_19_port, A2 => n1918, B1 => 
                           registers_30_19_port, B2 => n1915, ZN => n905);
   U1387 : AOI22_X1 port map( A1 => registers_23_20_port, A2 => n1941, B1 => 
                           registers_22_20_port, B2 => n1938, ZN => n920);
   U1388 : AOI22_X1 port map( A1 => registers_25_20_port, A2 => n1929, B1 => 
                           registers_24_20_port, B2 => n1926, ZN => n921);
   U1389 : AOI22_X1 port map( A1 => registers_31_20_port, A2 => n1917, B1 => 
                           registers_30_20_port, B2 => n1914, ZN => n922);
   U1390 : AOI22_X1 port map( A1 => registers_23_21_port, A2 => n1941, B1 => 
                           registers_22_21_port, B2 => n1938, ZN => n937);
   U1391 : AOI22_X1 port map( A1 => registers_25_21_port, A2 => n1929, B1 => 
                           registers_24_21_port, B2 => n1926, ZN => n938);
   U1392 : AOI22_X1 port map( A1 => registers_31_21_port, A2 => n1917, B1 => 
                           registers_30_21_port, B2 => n1914, ZN => n939);
   U1393 : AOI22_X1 port map( A1 => registers_23_22_port, A2 => n1941, B1 => 
                           registers_22_22_port, B2 => n1938, ZN => n954);
   U1394 : AOI22_X1 port map( A1 => registers_25_22_port, A2 => n1929, B1 => 
                           registers_24_22_port, B2 => n1926, ZN => n955);
   U1395 : AOI22_X1 port map( A1 => registers_31_22_port, A2 => n1917, B1 => 
                           registers_30_22_port, B2 => n1914, ZN => n956);
   U1396 : AOI22_X1 port map( A1 => registers_23_23_port, A2 => n1941, B1 => 
                           registers_22_23_port, B2 => n1938, ZN => n971);
   U1397 : AOI22_X1 port map( A1 => registers_25_23_port, A2 => n1929, B1 => 
                           registers_24_23_port, B2 => n1926, ZN => n972);
   U1398 : AOI22_X1 port map( A1 => registers_31_23_port, A2 => n1917, B1 => 
                           registers_30_23_port, B2 => n1914, ZN => n973);
   U1399 : AOI22_X1 port map( A1 => registers_23_24_port, A2 => n1941, B1 => 
                           registers_22_24_port, B2 => n1938, ZN => n988);
   U1400 : AOI22_X1 port map( A1 => registers_25_24_port, A2 => n1929, B1 => 
                           registers_24_24_port, B2 => n1926, ZN => n989);
   U1401 : AOI22_X1 port map( A1 => registers_31_24_port, A2 => n1917, B1 => 
                           registers_30_24_port, B2 => n1914, ZN => n990);
   U1402 : AOI22_X1 port map( A1 => registers_23_25_port, A2 => n1941, B1 => 
                           registers_22_25_port, B2 => n1938, ZN => n1005);
   U1403 : AOI22_X1 port map( A1 => registers_25_25_port, A2 => n1929, B1 => 
                           registers_24_25_port, B2 => n1926, ZN => n1006);
   U1404 : AOI22_X1 port map( A1 => registers_31_25_port, A2 => n1917, B1 => 
                           registers_30_25_port, B2 => n1914, ZN => n1007);
   U1405 : AOI22_X1 port map( A1 => registers_23_26_port, A2 => n1941, B1 => 
                           registers_22_26_port, B2 => n1938, ZN => n1022);
   U1406 : AOI22_X1 port map( A1 => registers_25_26_port, A2 => n1929, B1 => 
                           registers_24_26_port, B2 => n1926, ZN => n1023);
   U1407 : AOI22_X1 port map( A1 => registers_31_26_port, A2 => n1917, B1 => 
                           registers_30_26_port, B2 => n1914, ZN => n1024);
   U1408 : AOI22_X1 port map( A1 => registers_23_27_port, A2 => n1941, B1 => 
                           registers_22_27_port, B2 => n1938, ZN => n1039);
   U1409 : AOI22_X1 port map( A1 => registers_25_27_port, A2 => n1929, B1 => 
                           registers_24_27_port, B2 => n1926, ZN => n1040);
   U1410 : AOI22_X1 port map( A1 => registers_31_27_port, A2 => n1917, B1 => 
                           registers_30_27_port, B2 => n1914, ZN => n1041);
   U1411 : AOI22_X1 port map( A1 => registers_23_28_port, A2 => n1941, B1 => 
                           registers_22_28_port, B2 => n1938, ZN => n1056);
   U1412 : AOI22_X1 port map( A1 => registers_25_28_port, A2 => n1929, B1 => 
                           registers_24_28_port, B2 => n1926, ZN => n1057);
   U1413 : AOI22_X1 port map( A1 => registers_31_28_port, A2 => n1917, B1 => 
                           registers_30_28_port, B2 => n1914, ZN => n1058);
   U1414 : AOI22_X1 port map( A1 => registers_23_29_port, A2 => n1941, B1 => 
                           registers_22_29_port, B2 => n1938, ZN => n1073);
   U1415 : AOI22_X1 port map( A1 => registers_25_29_port, A2 => n1929, B1 => 
                           registers_24_29_port, B2 => n1926, ZN => n1074);
   U1416 : AOI22_X1 port map( A1 => registers_31_29_port, A2 => n1917, B1 => 
                           registers_30_29_port, B2 => n1914, ZN => n1075);
   U1417 : AOI22_X1 port map( A1 => registers_23_30_port, A2 => n1941, B1 => 
                           registers_22_30_port, B2 => n1938, ZN => n1090);
   U1418 : AOI22_X1 port map( A1 => registers_25_30_port, A2 => n1929, B1 => 
                           registers_24_30_port, B2 => n1926, ZN => n1091);
   U1419 : AOI22_X1 port map( A1 => registers_31_30_port, A2 => n1917, B1 => 
                           registers_30_30_port, B2 => n1914, ZN => n1092);
   U1420 : AOI22_X1 port map( A1 => registers_23_31_port, A2 => n1941, B1 => 
                           registers_22_31_port, B2 => n1938, ZN => n1111);
   U1421 : AOI22_X1 port map( A1 => registers_25_31_port, A2 => n1929, B1 => 
                           registers_24_31_port, B2 => n1926, ZN => n1114);
   U1422 : AOI22_X1 port map( A1 => registers_31_31_port, A2 => n1917, B1 => 
                           registers_30_31_port, B2 => n1914, ZN => n1117);
   U1423 : AND3_X1 port map( A1 => add_rd1(3), A2 => add_rd1(0), A3 => 
                           add_rd1(4), ZN => n1703);
   U1424 : AND3_X1 port map( A1 => add_rd1(3), A2 => n2684, A3 => add_rd1(4), 
                           ZN => n1702);
   U1425 : AND3_X1 port map( A1 => add_rd2(3), A2 => add_rd2(0), A3 => 
                           add_rd2(4), ZN => n1116);
   U1426 : AND3_X1 port map( A1 => n2684, A2 => n2681, A3 => add_rd1(4), ZN => 
                           n1694);
   U1427 : AND3_X1 port map( A1 => add_rd1(0), A2 => n2681, A3 => add_rd1(4), 
                           ZN => n1696);
   U1428 : AND3_X1 port map( A1 => add_rd2(3), A2 => n2688, A3 => add_rd2(4), 
                           ZN => n1115);
   U1429 : AND3_X1 port map( A1 => add_rd2(0), A2 => n2685, A3 => add_rd2(4), 
                           ZN => n1109);
   U1430 : AND3_X1 port map( A1 => n2688, A2 => n2685, A3 => add_rd2(4), ZN => 
                           n1107);
   U1431 : INV_X1 port map( A => add_rd2(3), ZN => n2685);
   U1432 : INV_X1 port map( A => add_rd2(0), ZN => n2688);
   U1433 : NAND4_X1 port map( A1 => n540, A2 => n541, A3 => n542, A4 => n543, 
                           ZN => N274);
   U1434 : AOI211_X1 port map( C1 => registers_5_0_port, C2 => n1913, A => n569
                           , B => n570, ZN => n542);
   U1435 : AOI221_X1 port map( B1 => registers_13_0_port, B2 => n1880, C1 => 
                           registers_2_0_port, C2 => n1877, A => n585, ZN => 
                           n540);
   U1436 : AOI221_X1 port map( B1 => registers_15_0_port, B2 => n1892, C1 => 
                           registers_12_0_port, C2 => n1889, A => n580, ZN => 
                           n541);
   U1437 : NAND4_X1 port map( A1 => n588, A2 => n589, A3 => n590, A4 => n591, 
                           ZN => N273);
   U1438 : AOI211_X1 port map( C1 => registers_5_1_port, C2 => n1913, A => n600
                           , B => n601, ZN => n590);
   U1439 : AOI221_X1 port map( B1 => registers_13_1_port, B2 => n1880, C1 => 
                           registers_2_1_port, C2 => n1877, A => n604, ZN => 
                           n588);
   U1440 : AOI221_X1 port map( B1 => registers_15_1_port, B2 => n1892, C1 => 
                           registers_12_1_port, C2 => n1889, A => n603, ZN => 
                           n589);
   U1441 : NAND4_X1 port map( A1 => n605, A2 => n606, A3 => n607, A4 => n608, 
                           ZN => N272);
   U1442 : AOI211_X1 port map( C1 => registers_5_2_port, C2 => n1913, A => n617
                           , B => n618, ZN => n607);
   U1443 : AOI221_X1 port map( B1 => registers_13_2_port, B2 => n1880, C1 => 
                           registers_2_2_port, C2 => n1877, A => n621, ZN => 
                           n605);
   U1444 : AOI221_X1 port map( B1 => registers_15_2_port, B2 => n1892, C1 => 
                           registers_12_2_port, C2 => n1889, A => n620, ZN => 
                           n606);
   U1445 : NAND4_X1 port map( A1 => n622, A2 => n623, A3 => n624, A4 => n625, 
                           ZN => N271);
   U1446 : AOI211_X1 port map( C1 => registers_5_3_port, C2 => n1913, A => n634
                           , B => n635, ZN => n624);
   U1447 : AOI221_X1 port map( B1 => registers_13_3_port, B2 => n1880, C1 => 
                           registers_2_3_port, C2 => n1877, A => n638, ZN => 
                           n622);
   U1448 : AOI221_X1 port map( B1 => registers_15_3_port, B2 => n1892, C1 => 
                           registers_12_3_port, C2 => n1889, A => n637, ZN => 
                           n623);
   U1449 : NAND4_X1 port map( A1 => n639, A2 => n640, A3 => n641, A4 => n642, 
                           ZN => N270);
   U1450 : AOI211_X1 port map( C1 => registers_5_4_port, C2 => n1913, A => n651
                           , B => n652, ZN => n641);
   U1451 : AOI221_X1 port map( B1 => registers_13_4_port, B2 => n1880, C1 => 
                           registers_2_4_port, C2 => n1877, A => n655, ZN => 
                           n639);
   U1452 : AOI221_X1 port map( B1 => registers_15_4_port, B2 => n1892, C1 => 
                           registers_12_4_port, C2 => n1889, A => n654, ZN => 
                           n640);
   U1453 : NAND4_X1 port map( A1 => n656, A2 => n657, A3 => n658, A4 => n659, 
                           ZN => N269);
   U1454 : AOI211_X1 port map( C1 => registers_5_5_port, C2 => n1913, A => n668
                           , B => n669, ZN => n658);
   U1455 : AOI221_X1 port map( B1 => registers_13_5_port, B2 => n1880, C1 => 
                           registers_2_5_port, C2 => n1877, A => n672, ZN => 
                           n656);
   U1456 : AOI221_X1 port map( B1 => registers_15_5_port, B2 => n1892, C1 => 
                           registers_12_5_port, C2 => n1889, A => n671, ZN => 
                           n657);
   U1457 : NAND4_X1 port map( A1 => n673, A2 => n674, A3 => n675, A4 => n676, 
                           ZN => N268);
   U1458 : AOI211_X1 port map( C1 => registers_5_6_port, C2 => n1913, A => n685
                           , B => n686, ZN => n675);
   U1459 : AOI221_X1 port map( B1 => registers_13_6_port, B2 => n1880, C1 => 
                           registers_2_6_port, C2 => n1877, A => n689, ZN => 
                           n673);
   U1460 : AOI221_X1 port map( B1 => registers_15_6_port, B2 => n1892, C1 => 
                           registers_12_6_port, C2 => n1889, A => n688, ZN => 
                           n674);
   U1461 : NAND4_X1 port map( A1 => n690, A2 => n691, A3 => n692, A4 => n693, 
                           ZN => N267);
   U1462 : AOI211_X1 port map( C1 => registers_5_7_port, C2 => n1913, A => n702
                           , B => n703, ZN => n692);
   U1463 : AOI221_X1 port map( B1 => registers_13_7_port, B2 => n1880, C1 => 
                           registers_2_7_port, C2 => n1877, A => n706, ZN => 
                           n690);
   U1464 : AOI221_X1 port map( B1 => registers_15_7_port, B2 => n1892, C1 => 
                           registers_12_7_port, C2 => n1889, A => n705, ZN => 
                           n691);
   U1465 : NAND4_X1 port map( A1 => n1127, A2 => n1128, A3 => n1129, A4 => 
                           n1130, ZN => N177);
   U1466 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_0_port, A => 
                           n1156, B => n1157, ZN => n1129);
   U1467 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_0_port, C1 => 
                           n1784, C2 => registers_2_0_port, A => n1172, ZN => 
                           n1127);
   U1468 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_0_port, C1 => 
                           n1796, C2 => registers_12_0_port, A => n1167, ZN => 
                           n1128);
   U1469 : NAND4_X1 port map( A1 => n1175, A2 => n1176, A3 => n1177, A4 => 
                           n1178, ZN => N176);
   U1470 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_1_port, A => 
                           n1187, B => n1188, ZN => n1177);
   U1471 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_1_port, C1 => 
                           n1784, C2 => registers_2_1_port, A => n1191, ZN => 
                           n1175);
   U1472 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_1_port, C1 => 
                           n1796, C2 => registers_12_1_port, A => n1190, ZN => 
                           n1176);
   U1473 : NAND4_X1 port map( A1 => n1192, A2 => n1193, A3 => n1194, A4 => 
                           n1195, ZN => N175);
   U1474 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_2_port, A => 
                           n1204, B => n1205, ZN => n1194);
   U1475 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_2_port, C1 => 
                           n1784, C2 => registers_2_2_port, A => n1208, ZN => 
                           n1192);
   U1476 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_2_port, C1 => 
                           n1796, C2 => registers_12_2_port, A => n1207, ZN => 
                           n1193);
   U1477 : NAND4_X1 port map( A1 => n1209, A2 => n1210, A3 => n1211, A4 => 
                           n1212, ZN => N174);
   U1478 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_3_port, A => 
                           n1221, B => n1222, ZN => n1211);
   U1479 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_3_port, C1 => 
                           n1784, C2 => registers_2_3_port, A => n1225, ZN => 
                           n1209);
   U1480 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_3_port, C1 => 
                           n1796, C2 => registers_12_3_port, A => n1224, ZN => 
                           n1210);
   U1481 : NAND4_X1 port map( A1 => n1226, A2 => n1227, A3 => n1228, A4 => 
                           n1229, ZN => N173);
   U1482 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_4_port, A => 
                           n1238, B => n1239, ZN => n1228);
   U1483 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_4_port, C1 => 
                           n1784, C2 => registers_2_4_port, A => n1242, ZN => 
                           n1226);
   U1484 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_4_port, C1 => 
                           n1796, C2 => registers_12_4_port, A => n1241, ZN => 
                           n1227);
   U1485 : NAND4_X1 port map( A1 => n1243, A2 => n1244, A3 => n1245, A4 => 
                           n1246, ZN => N172);
   U1486 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_5_port, A => 
                           n1255, B => n1256, ZN => n1245);
   U1487 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_5_port, C1 => 
                           n1784, C2 => registers_2_5_port, A => n1259, ZN => 
                           n1243);
   U1488 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_5_port, C1 => 
                           n1796, C2 => registers_12_5_port, A => n1258, ZN => 
                           n1244);
   U1489 : NAND4_X1 port map( A1 => n1260, A2 => n1261, A3 => n1262, A4 => 
                           n1263, ZN => N171);
   U1490 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_6_port, A => 
                           n1272, B => n1273, ZN => n1262);
   U1491 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_6_port, C1 => 
                           n1784, C2 => registers_2_6_port, A => n1276, ZN => 
                           n1260);
   U1492 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_6_port, C1 => 
                           n1796, C2 => registers_12_6_port, A => n1275, ZN => 
                           n1261);
   U1493 : NAND4_X1 port map( A1 => n1277, A2 => n1278, A3 => n1279, A4 => 
                           n1280, ZN => N170);
   U1494 : AOI211_X1 port map( C1 => n1820, C2 => registers_5_7_port, A => 
                           n1289, B => n1290, ZN => n1279);
   U1495 : AOI221_X1 port map( B1 => n1787, B2 => registers_13_7_port, C1 => 
                           n1784, C2 => registers_2_7_port, A => n1293, ZN => 
                           n1277);
   U1496 : AOI221_X1 port map( B1 => n1799, B2 => registers_15_7_port, C1 => 
                           n1796, C2 => registers_12_7_port, A => n1292, ZN => 
                           n1278);
   U1497 : NAND4_X1 port map( A1 => n1294, A2 => n1295, A3 => n1296, A4 => 
                           n1297, ZN => N169);
   U1498 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_8_port, A => 
                           n1306, B => n1307, ZN => n1296);
   U1499 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_8_port, C1 => 
                           n1783, C2 => registers_2_8_port, A => n1310, ZN => 
                           n1294);
   U1500 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_8_port, C1 => 
                           n1795, C2 => registers_12_8_port, A => n1309, ZN => 
                           n1295);
   U1501 : NAND4_X1 port map( A1 => n1311, A2 => n1312, A3 => n1313, A4 => 
                           n1314, ZN => N168);
   U1502 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_9_port, A => 
                           n1323, B => n1324, ZN => n1313);
   U1503 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_9_port, C1 => 
                           n1783, C2 => registers_2_9_port, A => n1327, ZN => 
                           n1311);
   U1504 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_9_port, C1 => 
                           n1795, C2 => registers_12_9_port, A => n1326, ZN => 
                           n1312);
   U1505 : NAND4_X1 port map( A1 => n1328, A2 => n1329, A3 => n1330, A4 => 
                           n1331, ZN => N167);
   U1506 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_10_port, A => 
                           n1340, B => n1341, ZN => n1330);
   U1507 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_10_port, C1 => 
                           n1783, C2 => registers_2_10_port, A => n1344, ZN => 
                           n1328);
   U1508 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_10_port, C1 => 
                           n1795, C2 => registers_12_10_port, A => n1343, ZN =>
                           n1329);
   U1509 : NAND4_X1 port map( A1 => n1345, A2 => n1346, A3 => n1347, A4 => 
                           n1348, ZN => N166);
   U1510 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_11_port, A => 
                           n1357, B => n1358, ZN => n1347);
   U1511 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_11_port, C1 => 
                           n1783, C2 => registers_2_11_port, A => n1361, ZN => 
                           n1345);
   U1512 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_11_port, C1 => 
                           n1795, C2 => registers_12_11_port, A => n1360, ZN =>
                           n1346);
   U1513 : NAND4_X1 port map( A1 => n1362, A2 => n1363, A3 => n1364, A4 => 
                           n1365, ZN => N165);
   U1514 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_12_port, A => 
                           n1374, B => n1375, ZN => n1364);
   U1515 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_12_port, C1 => 
                           n1783, C2 => registers_2_12_port, A => n1378, ZN => 
                           n1362);
   U1516 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_12_port, C1 => 
                           n1795, C2 => registers_12_12_port, A => n1377, ZN =>
                           n1363);
   U1517 : NAND4_X1 port map( A1 => n1379, A2 => n1380, A3 => n1381, A4 => 
                           n1382, ZN => N164);
   U1518 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_13_port, A => 
                           n1391, B => n1392, ZN => n1381);
   U1519 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_13_port, C1 => 
                           n1783, C2 => registers_2_13_port, A => n1395, ZN => 
                           n1379);
   U1520 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_13_port, C1 => 
                           n1795, C2 => registers_12_13_port, A => n1394, ZN =>
                           n1380);
   U1521 : NAND4_X1 port map( A1 => n1396, A2 => n1397, A3 => n1398, A4 => 
                           n1399, ZN => N163);
   U1522 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_14_port, A => 
                           n1408, B => n1409, ZN => n1398);
   U1523 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_14_port, C1 => 
                           n1783, C2 => registers_2_14_port, A => n1412, ZN => 
                           n1396);
   U1524 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_14_port, C1 => 
                           n1795, C2 => registers_12_14_port, A => n1411, ZN =>
                           n1397);
   U1525 : NAND4_X1 port map( A1 => n1413, A2 => n1414, A3 => n1415, A4 => 
                           n1416, ZN => N162);
   U1526 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_15_port, A => 
                           n1425, B => n1426, ZN => n1415);
   U1527 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_15_port, C1 => 
                           n1783, C2 => registers_2_15_port, A => n1429, ZN => 
                           n1413);
   U1528 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_15_port, C1 => 
                           n1795, C2 => registers_12_15_port, A => n1428, ZN =>
                           n1414);
   U1529 : NAND4_X1 port map( A1 => n1430, A2 => n1431, A3 => n1432, A4 => 
                           n1433, ZN => N161);
   U1530 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_16_port, A => 
                           n1442, B => n1443, ZN => n1432);
   U1531 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_16_port, C1 => 
                           n1783, C2 => registers_2_16_port, A => n1446, ZN => 
                           n1430);
   U1532 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_16_port, C1 => 
                           n1795, C2 => registers_12_16_port, A => n1445, ZN =>
                           n1431);
   U1533 : NAND4_X1 port map( A1 => n1447, A2 => n1448, A3 => n1449, A4 => 
                           n1450, ZN => N160);
   U1534 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_17_port, A => 
                           n1459, B => n1460, ZN => n1449);
   U1535 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_17_port, C1 => 
                           n1783, C2 => registers_2_17_port, A => n1463, ZN => 
                           n1447);
   U1536 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_17_port, C1 => 
                           n1795, C2 => registers_12_17_port, A => n1462, ZN =>
                           n1448);
   U1537 : NAND4_X1 port map( A1 => n1464, A2 => n1465, A3 => n1466, A4 => 
                           n1467, ZN => N159);
   U1538 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_18_port, A => 
                           n1476, B => n1477, ZN => n1466);
   U1539 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_18_port, C1 => 
                           n1783, C2 => registers_2_18_port, A => n1480, ZN => 
                           n1464);
   U1540 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_18_port, C1 => 
                           n1795, C2 => registers_12_18_port, A => n1479, ZN =>
                           n1465);
   U1541 : NAND4_X1 port map( A1 => n1481, A2 => n1482, A3 => n1483, A4 => 
                           n1484, ZN => N158);
   U1542 : AOI211_X1 port map( C1 => n1819, C2 => registers_5_19_port, A => 
                           n1493, B => n1494, ZN => n1483);
   U1543 : AOI221_X1 port map( B1 => n1786, B2 => registers_13_19_port, C1 => 
                           n1783, C2 => registers_2_19_port, A => n1497, ZN => 
                           n1481);
   U1544 : AOI221_X1 port map( B1 => n1798, B2 => registers_15_19_port, C1 => 
                           n1795, C2 => registers_12_19_port, A => n1496, ZN =>
                           n1482);
   U1545 : NAND4_X1 port map( A1 => n1498, A2 => n1499, A3 => n1500, A4 => 
                           n1501, ZN => N157);
   U1546 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_20_port, A => 
                           n1510, B => n1511, ZN => n1500);
   U1547 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_20_port, C1 => 
                           n1782, C2 => registers_2_20_port, A => n1514, ZN => 
                           n1498);
   U1548 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_20_port, C1 => 
                           n1794, C2 => registers_12_20_port, A => n1513, ZN =>
                           n1499);
   U1549 : NAND4_X1 port map( A1 => n1515, A2 => n1516, A3 => n1517, A4 => 
                           n1518, ZN => N156);
   U1550 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_21_port, A => 
                           n1527, B => n1528, ZN => n1517);
   U1551 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_21_port, C1 => 
                           n1782, C2 => registers_2_21_port, A => n1531, ZN => 
                           n1515);
   U1552 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_21_port, C1 => 
                           n1794, C2 => registers_12_21_port, A => n1530, ZN =>
                           n1516);
   U1553 : NAND4_X1 port map( A1 => n1532, A2 => n1533, A3 => n1534, A4 => 
                           n1535, ZN => N155);
   U1554 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_22_port, A => 
                           n1544, B => n1545, ZN => n1534);
   U1555 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_22_port, C1 => 
                           n1782, C2 => registers_2_22_port, A => n1548, ZN => 
                           n1532);
   U1556 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_22_port, C1 => 
                           n1794, C2 => registers_12_22_port, A => n1547, ZN =>
                           n1533);
   U1557 : NAND4_X1 port map( A1 => n1549, A2 => n1550, A3 => n1551, A4 => 
                           n1552, ZN => N154);
   U1558 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_23_port, A => 
                           n1561, B => n1562, ZN => n1551);
   U1559 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_23_port, C1 => 
                           n1782, C2 => registers_2_23_port, A => n1565, ZN => 
                           n1549);
   U1560 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_23_port, C1 => 
                           n1794, C2 => registers_12_23_port, A => n1564, ZN =>
                           n1550);
   U1561 : NAND4_X1 port map( A1 => n1566, A2 => n1567, A3 => n1568, A4 => 
                           n1569, ZN => N153);
   U1562 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_24_port, A => 
                           n1578, B => n1579, ZN => n1568);
   U1563 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_24_port, C1 => 
                           n1782, C2 => registers_2_24_port, A => n1582, ZN => 
                           n1566);
   U1564 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_24_port, C1 => 
                           n1794, C2 => registers_12_24_port, A => n1581, ZN =>
                           n1567);
   U1565 : NAND4_X1 port map( A1 => n1583, A2 => n1584, A3 => n1585, A4 => 
                           n1586, ZN => N152);
   U1566 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_25_port, A => 
                           n1595, B => n1596, ZN => n1585);
   U1567 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_25_port, C1 => 
                           n1782, C2 => registers_2_25_port, A => n1599, ZN => 
                           n1583);
   U1568 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_25_port, C1 => 
                           n1794, C2 => registers_12_25_port, A => n1598, ZN =>
                           n1584);
   U1569 : NAND4_X1 port map( A1 => n1600, A2 => n1601, A3 => n1602, A4 => 
                           n1603, ZN => N151);
   U1570 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_26_port, A => 
                           n1612, B => n1613, ZN => n1602);
   U1571 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_26_port, C1 => 
                           n1782, C2 => registers_2_26_port, A => n1616, ZN => 
                           n1600);
   U1572 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_26_port, C1 => 
                           n1794, C2 => registers_12_26_port, A => n1615, ZN =>
                           n1601);
   U1573 : NAND4_X1 port map( A1 => n1617, A2 => n1618, A3 => n1619, A4 => 
                           n1620, ZN => N150);
   U1574 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_27_port, A => 
                           n1629, B => n1630, ZN => n1619);
   U1575 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_27_port, C1 => 
                           n1782, C2 => registers_2_27_port, A => n1633, ZN => 
                           n1617);
   U1576 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_27_port, C1 => 
                           n1794, C2 => registers_12_27_port, A => n1632, ZN =>
                           n1618);
   U1577 : NAND4_X1 port map( A1 => n1634, A2 => n1635, A3 => n1636, A4 => 
                           n1637, ZN => N149);
   U1578 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_28_port, A => 
                           n1646, B => n1647, ZN => n1636);
   U1579 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_28_port, C1 => 
                           n1782, C2 => registers_2_28_port, A => n1650, ZN => 
                           n1634);
   U1580 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_28_port, C1 => 
                           n1794, C2 => registers_12_28_port, A => n1649, ZN =>
                           n1635);
   U1581 : NAND4_X1 port map( A1 => n1651, A2 => n1652, A3 => n1653, A4 => 
                           n1654, ZN => N148);
   U1582 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_29_port, A => 
                           n1663, B => n1664, ZN => n1653);
   U1583 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_29_port, C1 => 
                           n1782, C2 => registers_2_29_port, A => n1667, ZN => 
                           n1651);
   U1584 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_29_port, C1 => 
                           n1794, C2 => registers_12_29_port, A => n1666, ZN =>
                           n1652);
   U1585 : NAND4_X1 port map( A1 => n1668, A2 => n1669, A3 => n1670, A4 => 
                           n1671, ZN => N147);
   U1586 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_30_port, A => 
                           n1680, B => n1681, ZN => n1670);
   U1587 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_30_port, C1 => 
                           n1782, C2 => registers_2_30_port, A => n1684, ZN => 
                           n1668);
   U1588 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_30_port, C1 => 
                           n1794, C2 => registers_12_30_port, A => n1683, ZN =>
                           n1669);
   U1589 : NAND4_X1 port map( A1 => n1685, A2 => n1686, A3 => n1687, A4 => 
                           n1688, ZN => N146);
   U1590 : AOI211_X1 port map( C1 => n1818, C2 => registers_5_31_port, A => 
                           n1705, B => n1706, ZN => n1687);
   U1591 : AOI221_X1 port map( B1 => n1785, B2 => registers_13_31_port, C1 => 
                           n1782, C2 => registers_2_31_port, A => n1713, ZN => 
                           n1685);
   U1592 : AOI221_X1 port map( B1 => n1797, B2 => registers_15_31_port, C1 => 
                           n1794, C2 => registers_12_31_port, A => n1711, ZN =>
                           n1686);
   U1593 : NAND4_X1 port map( A1 => n707, A2 => n708, A3 => n709, A4 => n710, 
                           ZN => N266);
   U1594 : AOI211_X1 port map( C1 => registers_5_8_port, C2 => n1912, A => n719
                           , B => n720, ZN => n709);
   U1595 : AOI221_X1 port map( B1 => registers_13_8_port, B2 => n1879, C1 => 
                           registers_2_8_port, C2 => n1876, A => n723, ZN => 
                           n707);
   U1596 : AOI221_X1 port map( B1 => registers_15_8_port, B2 => n1891, C1 => 
                           registers_12_8_port, C2 => n1888, A => n722, ZN => 
                           n708);
   U1597 : NAND4_X1 port map( A1 => n724, A2 => n725, A3 => n726, A4 => n727, 
                           ZN => N265);
   U1598 : AOI211_X1 port map( C1 => registers_5_9_port, C2 => n1912, A => n736
                           , B => n737, ZN => n726);
   U1599 : AOI221_X1 port map( B1 => registers_13_9_port, B2 => n1879, C1 => 
                           registers_2_9_port, C2 => n1876, A => n740, ZN => 
                           n724);
   U1600 : AOI221_X1 port map( B1 => registers_15_9_port, B2 => n1891, C1 => 
                           registers_12_9_port, C2 => n1888, A => n739, ZN => 
                           n725);
   U1601 : NAND4_X1 port map( A1 => n741, A2 => n742, A3 => n743, A4 => n744, 
                           ZN => N264);
   U1602 : AOI211_X1 port map( C1 => registers_5_10_port, C2 => n1912, A => 
                           n753, B => n754, ZN => n743);
   U1603 : AOI221_X1 port map( B1 => registers_13_10_port, B2 => n1879, C1 => 
                           registers_2_10_port, C2 => n1876, A => n757, ZN => 
                           n741);
   U1604 : AOI221_X1 port map( B1 => registers_15_10_port, B2 => n1891, C1 => 
                           registers_12_10_port, C2 => n1888, A => n756, ZN => 
                           n742);
   U1605 : NAND4_X1 port map( A1 => n758, A2 => n759, A3 => n760, A4 => n761, 
                           ZN => N263);
   U1606 : AOI211_X1 port map( C1 => registers_5_11_port, C2 => n1912, A => 
                           n770, B => n771, ZN => n760);
   U1607 : AOI221_X1 port map( B1 => registers_13_11_port, B2 => n1879, C1 => 
                           registers_2_11_port, C2 => n1876, A => n774, ZN => 
                           n758);
   U1608 : AOI221_X1 port map( B1 => registers_15_11_port, B2 => n1891, C1 => 
                           registers_12_11_port, C2 => n1888, A => n773, ZN => 
                           n759);
   U1609 : NAND4_X1 port map( A1 => n775, A2 => n776, A3 => n777, A4 => n778, 
                           ZN => N262);
   U1610 : AOI211_X1 port map( C1 => registers_5_12_port, C2 => n1912, A => 
                           n787, B => n788, ZN => n777);
   U1611 : AOI221_X1 port map( B1 => registers_13_12_port, B2 => n1879, C1 => 
                           registers_2_12_port, C2 => n1876, A => n791, ZN => 
                           n775);
   U1612 : AOI221_X1 port map( B1 => registers_15_12_port, B2 => n1891, C1 => 
                           registers_12_12_port, C2 => n1888, A => n790, ZN => 
                           n776);
   U1613 : NAND4_X1 port map( A1 => n792, A2 => n793, A3 => n794, A4 => n795, 
                           ZN => N261);
   U1614 : AOI211_X1 port map( C1 => registers_5_13_port, C2 => n1912, A => 
                           n804, B => n805, ZN => n794);
   U1615 : AOI221_X1 port map( B1 => registers_13_13_port, B2 => n1879, C1 => 
                           registers_2_13_port, C2 => n1876, A => n808, ZN => 
                           n792);
   U1616 : AOI221_X1 port map( B1 => registers_15_13_port, B2 => n1891, C1 => 
                           registers_12_13_port, C2 => n1888, A => n807, ZN => 
                           n793);
   U1617 : NAND4_X1 port map( A1 => n809, A2 => n810, A3 => n811, A4 => n812, 
                           ZN => N260);
   U1618 : AOI211_X1 port map( C1 => registers_5_14_port, C2 => n1912, A => 
                           n821, B => n822, ZN => n811);
   U1619 : AOI221_X1 port map( B1 => registers_13_14_port, B2 => n1879, C1 => 
                           registers_2_14_port, C2 => n1876, A => n825, ZN => 
                           n809);
   U1620 : AOI221_X1 port map( B1 => registers_15_14_port, B2 => n1891, C1 => 
                           registers_12_14_port, C2 => n1888, A => n824, ZN => 
                           n810);
   U1621 : NAND4_X1 port map( A1 => n826, A2 => n827, A3 => n828, A4 => n829, 
                           ZN => N259);
   U1622 : AOI211_X1 port map( C1 => registers_5_15_port, C2 => n1912, A => 
                           n838, B => n839, ZN => n828);
   U1623 : AOI221_X1 port map( B1 => registers_13_15_port, B2 => n1879, C1 => 
                           registers_2_15_port, C2 => n1876, A => n842, ZN => 
                           n826);
   U1624 : AOI221_X1 port map( B1 => registers_15_15_port, B2 => n1891, C1 => 
                           registers_12_15_port, C2 => n1888, A => n841, ZN => 
                           n827);
   U1625 : NAND4_X1 port map( A1 => n843, A2 => n844, A3 => n845, A4 => n846, 
                           ZN => N258);
   U1626 : AOI211_X1 port map( C1 => registers_5_16_port, C2 => n1912, A => 
                           n855, B => n856, ZN => n845);
   U1627 : AOI221_X1 port map( B1 => registers_13_16_port, B2 => n1879, C1 => 
                           registers_2_16_port, C2 => n1876, A => n859, ZN => 
                           n843);
   U1628 : AOI221_X1 port map( B1 => registers_15_16_port, B2 => n1891, C1 => 
                           registers_12_16_port, C2 => n1888, A => n858, ZN => 
                           n844);
   U1629 : NAND4_X1 port map( A1 => n860, A2 => n861, A3 => n862, A4 => n863, 
                           ZN => N257);
   U1630 : AOI211_X1 port map( C1 => registers_5_17_port, C2 => n1912, A => 
                           n872, B => n873, ZN => n862);
   U1631 : AOI221_X1 port map( B1 => registers_13_17_port, B2 => n1879, C1 => 
                           registers_2_17_port, C2 => n1876, A => n876, ZN => 
                           n860);
   U1632 : AOI221_X1 port map( B1 => registers_15_17_port, B2 => n1891, C1 => 
                           registers_12_17_port, C2 => n1888, A => n875, ZN => 
                           n861);
   U1633 : NAND4_X1 port map( A1 => n877, A2 => n878, A3 => n879, A4 => n880, 
                           ZN => N256);
   U1634 : AOI211_X1 port map( C1 => registers_5_18_port, C2 => n1912, A => 
                           n889, B => n890, ZN => n879);
   U1635 : AOI221_X1 port map( B1 => registers_13_18_port, B2 => n1879, C1 => 
                           registers_2_18_port, C2 => n1876, A => n893, ZN => 
                           n877);
   U1636 : AOI221_X1 port map( B1 => registers_15_18_port, B2 => n1891, C1 => 
                           registers_12_18_port, C2 => n1888, A => n892, ZN => 
                           n878);
   U1637 : NAND4_X1 port map( A1 => n894, A2 => n895, A3 => n896, A4 => n897, 
                           ZN => N255);
   U1638 : AOI211_X1 port map( C1 => registers_5_19_port, C2 => n1912, A => 
                           n906, B => n907, ZN => n896);
   U1639 : AOI221_X1 port map( B1 => registers_13_19_port, B2 => n1879, C1 => 
                           registers_2_19_port, C2 => n1876, A => n910, ZN => 
                           n894);
   U1640 : AOI221_X1 port map( B1 => registers_15_19_port, B2 => n1891, C1 => 
                           registers_12_19_port, C2 => n1888, A => n909, ZN => 
                           n895);
   U1641 : NAND4_X1 port map( A1 => n911, A2 => n912, A3 => n913, A4 => n914, 
                           ZN => N254);
   U1642 : AOI211_X1 port map( C1 => registers_5_20_port, C2 => n1911, A => 
                           n923, B => n924, ZN => n913);
   U1643 : AOI221_X1 port map( B1 => registers_13_20_port, B2 => n1878, C1 => 
                           registers_2_20_port, C2 => n1875, A => n927, ZN => 
                           n911);
   U1644 : AOI221_X1 port map( B1 => registers_15_20_port, B2 => n1890, C1 => 
                           registers_12_20_port, C2 => n1887, A => n926, ZN => 
                           n912);
   U1645 : NAND4_X1 port map( A1 => n928, A2 => n929, A3 => n930, A4 => n931, 
                           ZN => N253);
   U1646 : AOI211_X1 port map( C1 => registers_5_21_port, C2 => n1911, A => 
                           n940, B => n941, ZN => n930);
   U1647 : AOI221_X1 port map( B1 => registers_13_21_port, B2 => n1878, C1 => 
                           registers_2_21_port, C2 => n1875, A => n944, ZN => 
                           n928);
   U1648 : AOI221_X1 port map( B1 => registers_15_21_port, B2 => n1890, C1 => 
                           registers_12_21_port, C2 => n1887, A => n943, ZN => 
                           n929);
   U1649 : NAND4_X1 port map( A1 => n945, A2 => n946, A3 => n947, A4 => n948, 
                           ZN => N252);
   U1650 : AOI211_X1 port map( C1 => registers_5_22_port, C2 => n1911, A => 
                           n957, B => n958, ZN => n947);
   U1651 : AOI221_X1 port map( B1 => registers_13_22_port, B2 => n1878, C1 => 
                           registers_2_22_port, C2 => n1875, A => n961, ZN => 
                           n945);
   U1652 : AOI221_X1 port map( B1 => registers_15_22_port, B2 => n1890, C1 => 
                           registers_12_22_port, C2 => n1887, A => n960, ZN => 
                           n946);
   U1653 : NAND4_X1 port map( A1 => n962, A2 => n963, A3 => n964, A4 => n965, 
                           ZN => N251);
   U1654 : AOI211_X1 port map( C1 => registers_5_23_port, C2 => n1911, A => 
                           n974, B => n975, ZN => n964);
   U1655 : AOI221_X1 port map( B1 => registers_13_23_port, B2 => n1878, C1 => 
                           registers_2_23_port, C2 => n1875, A => n978, ZN => 
                           n962);
   U1656 : AOI221_X1 port map( B1 => registers_15_23_port, B2 => n1890, C1 => 
                           registers_12_23_port, C2 => n1887, A => n977, ZN => 
                           n963);
   U1657 : NAND4_X1 port map( A1 => n979, A2 => n980, A3 => n981, A4 => n982, 
                           ZN => N250);
   U1658 : AOI211_X1 port map( C1 => registers_5_24_port, C2 => n1911, A => 
                           n991, B => n992, ZN => n981);
   U1659 : AOI221_X1 port map( B1 => registers_13_24_port, B2 => n1878, C1 => 
                           registers_2_24_port, C2 => n1875, A => n995, ZN => 
                           n979);
   U1660 : AOI221_X1 port map( B1 => registers_15_24_port, B2 => n1890, C1 => 
                           registers_12_24_port, C2 => n1887, A => n994, ZN => 
                           n980);
   U1661 : NAND4_X1 port map( A1 => n996, A2 => n997, A3 => n998, A4 => n999, 
                           ZN => N249);
   U1662 : AOI211_X1 port map( C1 => registers_5_25_port, C2 => n1911, A => 
                           n1008, B => n1009, ZN => n998);
   U1663 : AOI221_X1 port map( B1 => registers_13_25_port, B2 => n1878, C1 => 
                           registers_2_25_port, C2 => n1875, A => n1012, ZN => 
                           n996);
   U1664 : AOI221_X1 port map( B1 => registers_15_25_port, B2 => n1890, C1 => 
                           registers_12_25_port, C2 => n1887, A => n1011, ZN =>
                           n997);
   U1665 : NAND4_X1 port map( A1 => n1013, A2 => n1014, A3 => n1015, A4 => 
                           n1016, ZN => N248);
   U1666 : AOI211_X1 port map( C1 => registers_5_26_port, C2 => n1911, A => 
                           n1025, B => n1026, ZN => n1015);
   U1667 : AOI221_X1 port map( B1 => registers_13_26_port, B2 => n1878, C1 => 
                           registers_2_26_port, C2 => n1875, A => n1029, ZN => 
                           n1013);
   U1668 : AOI221_X1 port map( B1 => registers_15_26_port, B2 => n1890, C1 => 
                           registers_12_26_port, C2 => n1887, A => n1028, ZN =>
                           n1014);
   U1669 : NAND4_X1 port map( A1 => n1030, A2 => n1031, A3 => n1032, A4 => 
                           n1033, ZN => N247);
   U1670 : AOI211_X1 port map( C1 => registers_5_27_port, C2 => n1911, A => 
                           n1042, B => n1043, ZN => n1032);
   U1671 : AOI221_X1 port map( B1 => registers_13_27_port, B2 => n1878, C1 => 
                           registers_2_27_port, C2 => n1875, A => n1046, ZN => 
                           n1030);
   U1672 : AOI221_X1 port map( B1 => registers_15_27_port, B2 => n1890, C1 => 
                           registers_12_27_port, C2 => n1887, A => n1045, ZN =>
                           n1031);
   U1673 : NAND4_X1 port map( A1 => n1047, A2 => n1048, A3 => n1049, A4 => 
                           n1050, ZN => N246);
   U1674 : AOI211_X1 port map( C1 => registers_5_28_port, C2 => n1911, A => 
                           n1059, B => n1060, ZN => n1049);
   U1675 : AOI221_X1 port map( B1 => registers_13_28_port, B2 => n1878, C1 => 
                           registers_2_28_port, C2 => n1875, A => n1063, ZN => 
                           n1047);
   U1676 : AOI221_X1 port map( B1 => registers_15_28_port, B2 => n1890, C1 => 
                           registers_12_28_port, C2 => n1887, A => n1062, ZN =>
                           n1048);
   U1677 : NAND4_X1 port map( A1 => n1064, A2 => n1065, A3 => n1066, A4 => 
                           n1067, ZN => N245);
   U1678 : AOI211_X1 port map( C1 => registers_5_29_port, C2 => n1911, A => 
                           n1076, B => n1077, ZN => n1066);
   U1679 : AOI221_X1 port map( B1 => registers_13_29_port, B2 => n1878, C1 => 
                           registers_2_29_port, C2 => n1875, A => n1080, ZN => 
                           n1064);
   U1680 : AOI221_X1 port map( B1 => registers_15_29_port, B2 => n1890, C1 => 
                           registers_12_29_port, C2 => n1887, A => n1079, ZN =>
                           n1065);
   U1681 : NAND4_X1 port map( A1 => n1081, A2 => n1082, A3 => n1083, A4 => 
                           n1084, ZN => N244);
   U1682 : AOI211_X1 port map( C1 => registers_5_30_port, C2 => n1911, A => 
                           n1093, B => n1094, ZN => n1083);
   U1683 : AOI221_X1 port map( B1 => registers_13_30_port, B2 => n1878, C1 => 
                           registers_2_30_port, C2 => n1875, A => n1097, ZN => 
                           n1081);
   U1684 : AOI221_X1 port map( B1 => registers_15_30_port, B2 => n1890, C1 => 
                           registers_12_30_port, C2 => n1887, A => n1096, ZN =>
                           n1082);
   U1685 : NAND4_X1 port map( A1 => n1098, A2 => n1099, A3 => n1100, A4 => 
                           n1101, ZN => N243);
   U1686 : AOI211_X1 port map( C1 => registers_5_31_port, C2 => n1911, A => 
                           n1118, B => n1119, ZN => n1100);
   U1687 : AOI221_X1 port map( B1 => registers_13_31_port, B2 => n1878, C1 => 
                           registers_2_31_port, C2 => n1875, A => n1126, ZN => 
                           n1098);
   U1688 : AOI221_X1 port map( B1 => registers_15_31_port, B2 => n1890, C1 => 
                           registers_12_31_port, C2 => n1887, A => n1124, ZN =>
                           n1099);
   U1689 : INV_X1 port map( A => add_rd1(3), ZN => n2681);
   U1690 : INV_X1 port map( A => add_rd1(0), ZN => n2684);
   U1691 : INV_X1 port map( A => add_rd2(2), ZN => n2686);
   U1692 : INV_X1 port map( A => add_rd2(1), ZN => n2687);
   U1693 : INV_X1 port map( A => add_wr(2), ZN => n2166);
   U1694 : INV_X1 port map( A => add_wr(0), ZN => n2168);
   U1695 : INV_X1 port map( A => add_wr(1), ZN => n2167);
   U1696 : INV_X1 port map( A => add_rd1(2), ZN => n2682);
   U1697 : INV_X1 port map( A => add_rd1(1), ZN => n2683);
   U1698 : INV_X1 port map( A => registers_19_0_port, ZN => n2488);
   U1699 : INV_X1 port map( A => registers_21_0_port, ZN => n2552);
   U1700 : INV_X1 port map( A => registers_27_0_port, ZN => n2616);
   U1701 : INV_X1 port map( A => registers_29_0_port, ZN => n2680);
   U1702 : INV_X1 port map( A => registers_1_0_port, ZN => n2200);
   U1703 : INV_X1 port map( A => registers_19_1_port, ZN => n2487);
   U1704 : INV_X1 port map( A => registers_21_1_port, ZN => n2551);
   U1705 : INV_X1 port map( A => registers_27_1_port, ZN => n2615);
   U1706 : INV_X1 port map( A => registers_29_1_port, ZN => n2679);
   U1707 : INV_X1 port map( A => registers_1_1_port, ZN => n2199);
   U1708 : INV_X1 port map( A => registers_19_2_port, ZN => n2486);
   U1709 : INV_X1 port map( A => registers_21_2_port, ZN => n2550);
   U1710 : INV_X1 port map( A => registers_27_2_port, ZN => n2614);
   U1711 : INV_X1 port map( A => registers_29_2_port, ZN => n2678);
   U1712 : INV_X1 port map( A => registers_1_2_port, ZN => n2198);
   U1713 : INV_X1 port map( A => registers_19_3_port, ZN => n2485);
   U1714 : INV_X1 port map( A => registers_21_3_port, ZN => n2549);
   U1715 : INV_X1 port map( A => registers_27_3_port, ZN => n2613);
   U1716 : INV_X1 port map( A => registers_29_3_port, ZN => n2677);
   U1717 : INV_X1 port map( A => registers_1_3_port, ZN => n2197);
   U1718 : INV_X1 port map( A => registers_19_4_port, ZN => n2484);
   U1719 : INV_X1 port map( A => registers_21_4_port, ZN => n2548);
   U1720 : INV_X1 port map( A => registers_27_4_port, ZN => n2612);
   U1721 : INV_X1 port map( A => registers_29_4_port, ZN => n2676);
   U1722 : INV_X1 port map( A => registers_1_4_port, ZN => n2196);
   U1723 : INV_X1 port map( A => registers_19_5_port, ZN => n2483);
   U1724 : INV_X1 port map( A => registers_21_5_port, ZN => n2547);
   U1725 : INV_X1 port map( A => registers_27_5_port, ZN => n2611);
   U1726 : INV_X1 port map( A => registers_29_5_port, ZN => n2675);
   U1727 : INV_X1 port map( A => registers_1_5_port, ZN => n2195);
   U1728 : INV_X1 port map( A => registers_19_6_port, ZN => n2482);
   U1729 : INV_X1 port map( A => registers_21_6_port, ZN => n2546);
   U1730 : INV_X1 port map( A => registers_27_6_port, ZN => n2610);
   U1731 : INV_X1 port map( A => registers_29_6_port, ZN => n2674);
   U1732 : INV_X1 port map( A => registers_1_6_port, ZN => n2194);
   U1733 : INV_X1 port map( A => registers_19_7_port, ZN => n2481);
   U1734 : INV_X1 port map( A => registers_21_7_port, ZN => n2545);
   U1735 : INV_X1 port map( A => registers_27_7_port, ZN => n2609);
   U1736 : INV_X1 port map( A => registers_29_7_port, ZN => n2673);
   U1737 : INV_X1 port map( A => registers_1_7_port, ZN => n2193);
   U1738 : INV_X1 port map( A => registers_19_8_port, ZN => n2480);
   U1739 : INV_X1 port map( A => registers_21_8_port, ZN => n2544);
   U1740 : INV_X1 port map( A => registers_27_8_port, ZN => n2608);
   U1741 : INV_X1 port map( A => registers_29_8_port, ZN => n2672);
   U1742 : INV_X1 port map( A => registers_1_8_port, ZN => n2192);
   U1743 : INV_X1 port map( A => registers_19_9_port, ZN => n2479);
   U1744 : INV_X1 port map( A => registers_21_9_port, ZN => n2543);
   U1745 : INV_X1 port map( A => registers_27_9_port, ZN => n2607);
   U1746 : INV_X1 port map( A => registers_29_9_port, ZN => n2671);
   U1747 : INV_X1 port map( A => registers_1_9_port, ZN => n2191);
   U1748 : INV_X1 port map( A => registers_19_10_port, ZN => n2478);
   U1749 : INV_X1 port map( A => registers_21_10_port, ZN => n2542);
   U1750 : INV_X1 port map( A => registers_27_10_port, ZN => n2606);
   U1751 : INV_X1 port map( A => registers_29_10_port, ZN => n2670);
   U1752 : INV_X1 port map( A => registers_1_10_port, ZN => n2190);
   U1753 : INV_X1 port map( A => registers_19_11_port, ZN => n2477);
   U1754 : INV_X1 port map( A => registers_21_11_port, ZN => n2541);
   U1755 : INV_X1 port map( A => registers_27_11_port, ZN => n2605);
   U1756 : INV_X1 port map( A => registers_29_11_port, ZN => n2669);
   U1757 : INV_X1 port map( A => registers_1_11_port, ZN => n2189);
   U1758 : INV_X1 port map( A => registers_19_12_port, ZN => n2476);
   U1759 : INV_X1 port map( A => registers_21_12_port, ZN => n2540);
   U1760 : INV_X1 port map( A => registers_27_12_port, ZN => n2604);
   U1761 : INV_X1 port map( A => registers_29_12_port, ZN => n2668);
   U1762 : INV_X1 port map( A => registers_1_12_port, ZN => n2188);
   U1763 : INV_X1 port map( A => registers_19_13_port, ZN => n2475);
   U1764 : INV_X1 port map( A => registers_21_13_port, ZN => n2539);
   U1765 : INV_X1 port map( A => registers_27_13_port, ZN => n2603);
   U1766 : INV_X1 port map( A => registers_29_13_port, ZN => n2667);
   U1767 : INV_X1 port map( A => registers_1_13_port, ZN => n2187);
   U1768 : INV_X1 port map( A => registers_19_14_port, ZN => n2474);
   U1769 : INV_X1 port map( A => registers_21_14_port, ZN => n2538);
   U1770 : INV_X1 port map( A => registers_27_14_port, ZN => n2602);
   U1771 : INV_X1 port map( A => registers_29_14_port, ZN => n2666);
   U1772 : INV_X1 port map( A => registers_1_14_port, ZN => n2186);
   U1773 : INV_X1 port map( A => registers_19_15_port, ZN => n2473);
   U1774 : INV_X1 port map( A => registers_21_15_port, ZN => n2537);
   U1775 : INV_X1 port map( A => registers_27_15_port, ZN => n2601);
   U1776 : INV_X1 port map( A => registers_29_15_port, ZN => n2665);
   U1777 : INV_X1 port map( A => registers_1_15_port, ZN => n2185);
   U1778 : INV_X1 port map( A => registers_19_16_port, ZN => n2472);
   U1779 : INV_X1 port map( A => registers_21_16_port, ZN => n2536);
   U1780 : INV_X1 port map( A => registers_27_16_port, ZN => n2600);
   U1781 : INV_X1 port map( A => registers_29_16_port, ZN => n2664);
   U1782 : INV_X1 port map( A => registers_1_16_port, ZN => n2184);
   U1783 : INV_X1 port map( A => registers_19_17_port, ZN => n2471);
   U1784 : INV_X1 port map( A => registers_21_17_port, ZN => n2535);
   U1785 : INV_X1 port map( A => registers_27_17_port, ZN => n2599);
   U1786 : INV_X1 port map( A => registers_29_17_port, ZN => n2663);
   U1787 : INV_X1 port map( A => registers_1_17_port, ZN => n2183);
   U1788 : INV_X1 port map( A => registers_19_18_port, ZN => n2470);
   U1789 : INV_X1 port map( A => registers_21_18_port, ZN => n2534);
   U1790 : INV_X1 port map( A => registers_27_18_port, ZN => n2598);
   U1791 : INV_X1 port map( A => registers_29_18_port, ZN => n2662);
   U1792 : INV_X1 port map( A => registers_1_18_port, ZN => n2182);
   U1793 : INV_X1 port map( A => registers_19_19_port, ZN => n2469);
   U1794 : INV_X1 port map( A => registers_21_19_port, ZN => n2533);
   U1795 : INV_X1 port map( A => registers_27_19_port, ZN => n2597);
   U1796 : INV_X1 port map( A => registers_29_19_port, ZN => n2661);
   U1797 : INV_X1 port map( A => registers_1_19_port, ZN => n2181);
   U1798 : INV_X1 port map( A => registers_19_20_port, ZN => n2468);
   U1799 : INV_X1 port map( A => registers_21_20_port, ZN => n2532);
   U1800 : INV_X1 port map( A => registers_27_20_port, ZN => n2596);
   U1801 : INV_X1 port map( A => registers_29_20_port, ZN => n2660);
   U1802 : INV_X1 port map( A => registers_1_20_port, ZN => n2180);
   U1803 : INV_X1 port map( A => registers_19_21_port, ZN => n2467);
   U1804 : INV_X1 port map( A => registers_21_21_port, ZN => n2531);
   U1805 : INV_X1 port map( A => registers_27_21_port, ZN => n2595);
   U1806 : INV_X1 port map( A => registers_29_21_port, ZN => n2659);
   U1807 : INV_X1 port map( A => registers_1_21_port, ZN => n2179);
   U1808 : INV_X1 port map( A => registers_19_22_port, ZN => n2466);
   U1809 : INV_X1 port map( A => registers_21_22_port, ZN => n2530);
   U1810 : INV_X1 port map( A => registers_27_22_port, ZN => n2594);
   U1811 : INV_X1 port map( A => registers_29_22_port, ZN => n2658);
   U1812 : INV_X1 port map( A => registers_1_22_port, ZN => n2178);
   U1813 : INV_X1 port map( A => registers_19_23_port, ZN => n2465);
   U1814 : INV_X1 port map( A => registers_21_23_port, ZN => n2529);
   U1815 : INV_X1 port map( A => registers_27_23_port, ZN => n2593);
   U1816 : INV_X1 port map( A => registers_29_23_port, ZN => n2657);
   U1817 : INV_X1 port map( A => registers_1_23_port, ZN => n2177);
   U1818 : INV_X1 port map( A => registers_19_24_port, ZN => n2464);
   U1819 : INV_X1 port map( A => registers_21_24_port, ZN => n2528);
   U1820 : INV_X1 port map( A => registers_27_24_port, ZN => n2592);
   U1821 : INV_X1 port map( A => registers_29_24_port, ZN => n2656);
   U1822 : INV_X1 port map( A => registers_1_24_port, ZN => n2176);
   U1823 : INV_X1 port map( A => registers_19_25_port, ZN => n2463);
   U1824 : INV_X1 port map( A => registers_21_25_port, ZN => n2527);
   U1825 : INV_X1 port map( A => registers_27_25_port, ZN => n2591);
   U1826 : INV_X1 port map( A => registers_29_25_port, ZN => n2655);
   U1827 : INV_X1 port map( A => registers_1_25_port, ZN => n2175);
   U1828 : INV_X1 port map( A => registers_19_26_port, ZN => n2462);
   U1829 : INV_X1 port map( A => registers_21_26_port, ZN => n2526);
   U1830 : INV_X1 port map( A => registers_27_26_port, ZN => n2590);
   U1831 : INV_X1 port map( A => registers_29_26_port, ZN => n2654);
   U1844 : INV_X1 port map( A => registers_1_26_port, ZN => n2174);
   U1845 : INV_X1 port map( A => registers_19_27_port, ZN => n2461);
   U1846 : INV_X1 port map( A => registers_21_27_port, ZN => n2525);
   U1847 : INV_X1 port map( A => registers_27_27_port, ZN => n2589);
   U1848 : INV_X1 port map( A => registers_29_27_port, ZN => n2653);
   U1849 : INV_X1 port map( A => registers_1_27_port, ZN => n2173);
   U1850 : INV_X1 port map( A => registers_19_28_port, ZN => n2460);
   U1851 : INV_X1 port map( A => registers_21_28_port, ZN => n2524);
   U1852 : INV_X1 port map( A => registers_27_28_port, ZN => n2588);
   U1853 : INV_X1 port map( A => registers_29_28_port, ZN => n2652);
   U1854 : INV_X1 port map( A => registers_1_28_port, ZN => n2172);
   U1855 : INV_X1 port map( A => registers_19_29_port, ZN => n2459);
   U1856 : INV_X1 port map( A => registers_21_29_port, ZN => n2523);
   U1857 : INV_X1 port map( A => registers_27_29_port, ZN => n2587);
   U1858 : INV_X1 port map( A => registers_29_29_port, ZN => n2651);
   U1859 : INV_X1 port map( A => registers_1_29_port, ZN => n2171);
   U1860 : INV_X1 port map( A => registers_19_30_port, ZN => n2458);
   U1861 : INV_X1 port map( A => registers_21_30_port, ZN => n2522);
   U1862 : INV_X1 port map( A => registers_27_30_port, ZN => n2586);
   U1863 : INV_X1 port map( A => registers_29_30_port, ZN => n2650);
   U1864 : INV_X1 port map( A => registers_1_30_port, ZN => n2170);
   U1865 : INV_X1 port map( A => registers_19_31_port, ZN => n2457);
   U1866 : INV_X1 port map( A => registers_21_31_port, ZN => n2521);
   U1867 : INV_X1 port map( A => registers_27_31_port, ZN => n2585);
   U1868 : INV_X1 port map( A => registers_29_31_port, ZN => n2649);
   U1869 : INV_X1 port map( A => registers_1_31_port, ZN => n2169);
   U1870 : INV_X1 port map( A => registers_11_0_port, ZN => n2392);
   U1871 : INV_X1 port map( A => registers_9_0_port, ZN => n2328);
   U1872 : INV_X1 port map( A => registers_10_0_port, ZN => n2360);
   U1873 : INV_X1 port map( A => registers_11_1_port, ZN => n2391);
   U1874 : INV_X1 port map( A => registers_9_1_port, ZN => n2327);
   U1875 : INV_X1 port map( A => registers_10_1_port, ZN => n2359);
   U1876 : INV_X1 port map( A => registers_11_2_port, ZN => n2390);
   U1877 : INV_X1 port map( A => registers_9_2_port, ZN => n2326);
   U1878 : INV_X1 port map( A => registers_10_2_port, ZN => n2358);
   U1879 : INV_X1 port map( A => registers_11_3_port, ZN => n2389);
   U1880 : INV_X1 port map( A => registers_9_3_port, ZN => n2325);
   U1881 : INV_X1 port map( A => registers_10_3_port, ZN => n2357);
   U1882 : INV_X1 port map( A => registers_11_4_port, ZN => n2388);
   U1883 : INV_X1 port map( A => registers_9_4_port, ZN => n2324);
   U1884 : INV_X1 port map( A => registers_10_4_port, ZN => n2356);
   U1885 : INV_X1 port map( A => registers_11_5_port, ZN => n2387);
   U1886 : INV_X1 port map( A => registers_9_5_port, ZN => n2323);
   U1887 : INV_X1 port map( A => registers_10_5_port, ZN => n2355);
   U1888 : INV_X1 port map( A => registers_11_6_port, ZN => n2386);
   U1889 : INV_X1 port map( A => registers_9_6_port, ZN => n2322);
   U1890 : INV_X1 port map( A => registers_10_6_port, ZN => n2354);
   U1891 : INV_X1 port map( A => registers_11_7_port, ZN => n2385);
   U1892 : INV_X1 port map( A => registers_9_7_port, ZN => n2321);
   U1893 : INV_X1 port map( A => registers_10_7_port, ZN => n2353);
   U1894 : INV_X1 port map( A => registers_11_8_port, ZN => n2384);
   U1895 : INV_X1 port map( A => registers_9_8_port, ZN => n2320);
   U1896 : INV_X1 port map( A => registers_10_8_port, ZN => n2352);
   U1897 : INV_X1 port map( A => registers_11_9_port, ZN => n2383);
   U1898 : INV_X1 port map( A => registers_9_9_port, ZN => n2319);
   U1899 : INV_X1 port map( A => registers_10_9_port, ZN => n2351);
   U1900 : INV_X1 port map( A => registers_11_10_port, ZN => n2382);
   U1901 : INV_X1 port map( A => registers_9_10_port, ZN => n2318);
   U1902 : INV_X1 port map( A => registers_10_10_port, ZN => n2350);
   U1903 : INV_X1 port map( A => registers_11_11_port, ZN => n2381);
   U1904 : INV_X1 port map( A => registers_9_11_port, ZN => n2317);
   U1905 : INV_X1 port map( A => registers_10_11_port, ZN => n2349);
   U1906 : INV_X1 port map( A => registers_11_12_port, ZN => n2380);
   U1907 : INV_X1 port map( A => registers_9_12_port, ZN => n2316);
   U1908 : INV_X1 port map( A => registers_10_12_port, ZN => n2348);
   U1909 : INV_X1 port map( A => registers_11_13_port, ZN => n2379);
   U1910 : INV_X1 port map( A => registers_9_13_port, ZN => n2315);
   U1911 : INV_X1 port map( A => registers_10_13_port, ZN => n2347);
   U1912 : INV_X1 port map( A => registers_11_14_port, ZN => n2378);
   U1913 : INV_X1 port map( A => registers_9_14_port, ZN => n2314);
   U1914 : INV_X1 port map( A => registers_10_14_port, ZN => n2346);
   U1915 : INV_X1 port map( A => registers_11_15_port, ZN => n2377);
   U1916 : INV_X1 port map( A => registers_9_15_port, ZN => n2313);
   U1917 : INV_X1 port map( A => registers_10_15_port, ZN => n2345);
   U1918 : INV_X1 port map( A => registers_11_16_port, ZN => n2376);
   U1919 : INV_X1 port map( A => registers_9_16_port, ZN => n2312);
   U1920 : INV_X1 port map( A => registers_10_16_port, ZN => n2344);
   U1921 : INV_X1 port map( A => registers_11_17_port, ZN => n2375);
   U1922 : INV_X1 port map( A => registers_9_17_port, ZN => n2311);
   U1923 : INV_X1 port map( A => registers_10_17_port, ZN => n2343);
   U1924 : INV_X1 port map( A => registers_11_18_port, ZN => n2374);
   U1925 : INV_X1 port map( A => registers_9_18_port, ZN => n2310);
   U1926 : INV_X1 port map( A => registers_10_18_port, ZN => n2342);
   U1927 : INV_X1 port map( A => registers_11_19_port, ZN => n2373);
   U1928 : INV_X1 port map( A => registers_9_19_port, ZN => n2309);
   U1929 : INV_X1 port map( A => registers_10_19_port, ZN => n2341);
   U1930 : INV_X1 port map( A => registers_11_20_port, ZN => n2372);
   U1931 : INV_X1 port map( A => registers_9_20_port, ZN => n2308);
   U1932 : INV_X1 port map( A => registers_10_20_port, ZN => n2340);
   U1933 : INV_X1 port map( A => registers_11_21_port, ZN => n2371);
   U1934 : INV_X1 port map( A => registers_9_21_port, ZN => n2307);
   U1935 : INV_X1 port map( A => registers_10_21_port, ZN => n2339);
   U1936 : INV_X1 port map( A => registers_11_22_port, ZN => n2370);
   U1937 : INV_X1 port map( A => registers_9_22_port, ZN => n2306);
   U1938 : INV_X1 port map( A => registers_10_22_port, ZN => n2338);
   U1939 : INV_X1 port map( A => registers_11_23_port, ZN => n2369);
   U1940 : INV_X1 port map( A => registers_9_23_port, ZN => n2305);
   U1941 : INV_X1 port map( A => registers_10_23_port, ZN => n2337);
   U1942 : INV_X1 port map( A => registers_11_24_port, ZN => n2368);
   U1943 : INV_X1 port map( A => registers_9_24_port, ZN => n2304);
   U1944 : INV_X1 port map( A => registers_10_24_port, ZN => n2336);
   U1945 : INV_X1 port map( A => registers_11_25_port, ZN => n2367);
   U1946 : INV_X1 port map( A => registers_9_25_port, ZN => n2303);
   U1947 : INV_X1 port map( A => registers_10_25_port, ZN => n2335);
   U1948 : INV_X1 port map( A => registers_11_26_port, ZN => n2366);
   U1949 : INV_X1 port map( A => registers_9_26_port, ZN => n2302);
   U1950 : INV_X1 port map( A => registers_10_26_port, ZN => n2334);
   U1951 : INV_X1 port map( A => registers_11_27_port, ZN => n2365);
   U1952 : INV_X1 port map( A => registers_9_27_port, ZN => n2301);
   U1953 : INV_X1 port map( A => registers_10_27_port, ZN => n2333);
   U1954 : INV_X1 port map( A => registers_11_28_port, ZN => n2364);
   U1955 : INV_X1 port map( A => registers_9_28_port, ZN => n2300);
   U1956 : INV_X1 port map( A => registers_10_28_port, ZN => n2332);
   U1957 : INV_X1 port map( A => registers_11_29_port, ZN => n2363);
   U1958 : INV_X1 port map( A => registers_9_29_port, ZN => n2299);
   U1959 : INV_X1 port map( A => registers_10_29_port, ZN => n2331);
   U1960 : INV_X1 port map( A => registers_11_30_port, ZN => n2362);
   U1961 : INV_X1 port map( A => registers_9_30_port, ZN => n2298);
   U1962 : INV_X1 port map( A => registers_10_30_port, ZN => n2330);
   U1963 : INV_X1 port map( A => registers_11_31_port, ZN => n2361);
   U1964 : INV_X1 port map( A => registers_9_31_port, ZN => n2297);
   U1965 : INV_X1 port map( A => registers_10_31_port, ZN => n2329);
   U1966 : INV_X1 port map( A => registers_8_0_port, ZN => n2296);
   U1967 : INV_X1 port map( A => registers_14_0_port, ZN => n2424);
   U1968 : INV_X1 port map( A => registers_4_0_port, ZN => n2232);
   U1969 : INV_X1 port map( A => registers_8_1_port, ZN => n2295);
   U1970 : INV_X1 port map( A => registers_14_1_port, ZN => n2423);
   U1971 : INV_X1 port map( A => registers_4_1_port, ZN => n2231);
   U1972 : INV_X1 port map( A => registers_8_2_port, ZN => n2294);
   U1973 : INV_X1 port map( A => registers_14_2_port, ZN => n2422);
   U1974 : INV_X1 port map( A => registers_4_2_port, ZN => n2230);
   U1975 : INV_X1 port map( A => registers_8_3_port, ZN => n2293);
   U1976 : INV_X1 port map( A => registers_14_3_port, ZN => n2421);
   U1977 : INV_X1 port map( A => registers_4_3_port, ZN => n2229);
   U1978 : INV_X1 port map( A => registers_8_4_port, ZN => n2292);
   U1979 : INV_X1 port map( A => registers_14_4_port, ZN => n2420);
   U1980 : INV_X1 port map( A => registers_4_4_port, ZN => n2228);
   U1981 : INV_X1 port map( A => registers_8_5_port, ZN => n2291);
   U1982 : INV_X1 port map( A => registers_14_5_port, ZN => n2419);
   U1983 : INV_X1 port map( A => registers_4_5_port, ZN => n2227);
   U1984 : INV_X1 port map( A => registers_8_6_port, ZN => n2290);
   U1985 : INV_X1 port map( A => registers_14_6_port, ZN => n2418);
   U1986 : INV_X1 port map( A => registers_4_6_port, ZN => n2226);
   U1987 : INV_X1 port map( A => registers_8_7_port, ZN => n2289);
   U1988 : INV_X1 port map( A => registers_14_7_port, ZN => n2417);
   U1989 : INV_X1 port map( A => registers_4_7_port, ZN => n2225);
   U1990 : INV_X1 port map( A => registers_8_8_port, ZN => n2288);
   U1991 : INV_X1 port map( A => registers_14_8_port, ZN => n2416);
   U1992 : INV_X1 port map( A => registers_4_8_port, ZN => n2224);
   U1993 : INV_X1 port map( A => registers_8_9_port, ZN => n2287);
   U1994 : INV_X1 port map( A => registers_14_9_port, ZN => n2415);
   U1995 : INV_X1 port map( A => registers_4_9_port, ZN => n2223);
   U1996 : INV_X1 port map( A => registers_8_10_port, ZN => n2286);
   U1997 : INV_X1 port map( A => registers_14_10_port, ZN => n2414);
   U1998 : INV_X1 port map( A => registers_4_10_port, ZN => n2222);
   U1999 : INV_X1 port map( A => registers_8_11_port, ZN => n2285);
   U2000 : INV_X1 port map( A => registers_14_11_port, ZN => n2413);
   U2001 : INV_X1 port map( A => registers_4_11_port, ZN => n2221);
   U2002 : INV_X1 port map( A => registers_8_12_port, ZN => n2284);
   U2003 : INV_X1 port map( A => registers_14_12_port, ZN => n2412);
   U2004 : INV_X1 port map( A => registers_4_12_port, ZN => n2220);
   U2005 : INV_X1 port map( A => registers_8_13_port, ZN => n2283);
   U2006 : INV_X1 port map( A => registers_14_13_port, ZN => n2411);
   U2007 : INV_X1 port map( A => registers_4_13_port, ZN => n2219);
   U2008 : INV_X1 port map( A => registers_8_14_port, ZN => n2282);
   U2009 : INV_X1 port map( A => registers_14_14_port, ZN => n2410);
   U2010 : INV_X1 port map( A => registers_4_14_port, ZN => n2218);
   U2011 : INV_X1 port map( A => registers_8_15_port, ZN => n2281);
   U2012 : INV_X1 port map( A => registers_14_15_port, ZN => n2409);
   U2013 : INV_X1 port map( A => registers_4_15_port, ZN => n2217);
   U2014 : INV_X1 port map( A => registers_8_16_port, ZN => n2280);
   U2015 : INV_X1 port map( A => registers_14_16_port, ZN => n2408);
   U2016 : INV_X1 port map( A => registers_4_16_port, ZN => n2216);
   U2017 : INV_X1 port map( A => registers_8_17_port, ZN => n2279);
   U2018 : INV_X1 port map( A => registers_14_17_port, ZN => n2407);
   U2019 : INV_X1 port map( A => registers_4_17_port, ZN => n2215);
   U2020 : INV_X1 port map( A => registers_8_18_port, ZN => n2278);
   U2021 : INV_X1 port map( A => registers_14_18_port, ZN => n2406);
   U2022 : INV_X1 port map( A => registers_4_18_port, ZN => n2214);
   U2023 : INV_X1 port map( A => registers_8_19_port, ZN => n2277);
   U2024 : INV_X1 port map( A => registers_14_19_port, ZN => n2405);
   U2025 : INV_X1 port map( A => registers_4_19_port, ZN => n2213);
   U2026 : INV_X1 port map( A => registers_8_20_port, ZN => n2276);
   U2027 : INV_X1 port map( A => registers_14_20_port, ZN => n2404);
   U2028 : INV_X1 port map( A => registers_4_20_port, ZN => n2212);
   U2029 : INV_X1 port map( A => registers_8_21_port, ZN => n2275);
   U2030 : INV_X1 port map( A => registers_14_21_port, ZN => n2403);
   U2031 : INV_X1 port map( A => registers_4_21_port, ZN => n2211);
   U2032 : INV_X1 port map( A => registers_8_22_port, ZN => n2274);
   U2033 : INV_X1 port map( A => registers_14_22_port, ZN => n2402);
   U2034 : INV_X1 port map( A => registers_4_22_port, ZN => n2210);
   U2035 : INV_X1 port map( A => registers_8_23_port, ZN => n2273);
   U2036 : INV_X1 port map( A => registers_14_23_port, ZN => n2401);
   U2037 : INV_X1 port map( A => registers_4_23_port, ZN => n2209);
   U2038 : INV_X1 port map( A => registers_8_24_port, ZN => n2272);
   U2039 : INV_X1 port map( A => registers_14_24_port, ZN => n2400);
   U2040 : INV_X1 port map( A => registers_4_24_port, ZN => n2208);
   U2041 : INV_X1 port map( A => registers_8_25_port, ZN => n2271);
   U2042 : INV_X1 port map( A => registers_14_25_port, ZN => n2399);
   U2043 : INV_X1 port map( A => registers_4_25_port, ZN => n2207);
   U2044 : INV_X1 port map( A => registers_8_26_port, ZN => n2270);
   U2045 : INV_X1 port map( A => registers_14_26_port, ZN => n2398);
   U2046 : INV_X1 port map( A => registers_4_26_port, ZN => n2206);
   U2047 : INV_X1 port map( A => registers_8_27_port, ZN => n2269);
   U2048 : INV_X1 port map( A => registers_14_27_port, ZN => n2397);
   U2049 : INV_X1 port map( A => registers_4_27_port, ZN => n2205);
   U2050 : INV_X1 port map( A => registers_8_28_port, ZN => n2268);
   U2051 : INV_X1 port map( A => registers_14_28_port, ZN => n2396);
   U2052 : INV_X1 port map( A => registers_4_28_port, ZN => n2204);
   U2053 : INV_X1 port map( A => registers_8_29_port, ZN => n2267);
   U2054 : INV_X1 port map( A => registers_14_29_port, ZN => n2395);
   U2055 : INV_X1 port map( A => registers_4_29_port, ZN => n2203);
   U2056 : INV_X1 port map( A => registers_8_30_port, ZN => n2266);
   U2057 : INV_X1 port map( A => registers_14_30_port, ZN => n2394);
   U2058 : INV_X1 port map( A => registers_4_30_port, ZN => n2202);
   U2059 : INV_X1 port map( A => registers_8_31_port, ZN => n2265);
   U2060 : INV_X1 port map( A => registers_14_31_port, ZN => n2393);
   U2061 : INV_X1 port map( A => registers_4_31_port, ZN => n2201);
   U2062 : INV_X1 port map( A => registers_18_0_port, ZN => n2456);
   U2063 : INV_X1 port map( A => registers_20_0_port, ZN => n2520);
   U2064 : INV_X1 port map( A => registers_26_0_port, ZN => n2584);
   U2065 : INV_X1 port map( A => registers_28_0_port, ZN => n2648);
   U2066 : INV_X1 port map( A => registers_7_0_port, ZN => n2264);
   U2067 : INV_X1 port map( A => registers_18_1_port, ZN => n2455);
   U2068 : INV_X1 port map( A => registers_20_1_port, ZN => n2519);
   U2069 : INV_X1 port map( A => registers_26_1_port, ZN => n2583);
   U2070 : INV_X1 port map( A => registers_28_1_port, ZN => n2647);
   U2071 : INV_X1 port map( A => registers_7_1_port, ZN => n2263);
   U2072 : INV_X1 port map( A => registers_18_2_port, ZN => n2454);
   U2073 : INV_X1 port map( A => registers_20_2_port, ZN => n2518);
   U2074 : INV_X1 port map( A => registers_26_2_port, ZN => n2582);
   U2075 : INV_X1 port map( A => registers_28_2_port, ZN => n2646);
   U2076 : INV_X1 port map( A => registers_7_2_port, ZN => n2262);
   U2077 : INV_X1 port map( A => registers_18_3_port, ZN => n2453);
   U2078 : INV_X1 port map( A => registers_20_3_port, ZN => n2517);
   U2079 : INV_X1 port map( A => registers_26_3_port, ZN => n2581);
   U2080 : INV_X1 port map( A => registers_28_3_port, ZN => n2645);
   U2081 : INV_X1 port map( A => registers_7_3_port, ZN => n2261);
   U2082 : INV_X1 port map( A => registers_18_4_port, ZN => n2452);
   U2083 : INV_X1 port map( A => registers_20_4_port, ZN => n2516);
   U2084 : INV_X1 port map( A => registers_26_4_port, ZN => n2580);
   U2085 : INV_X1 port map( A => registers_28_4_port, ZN => n2644);
   U2086 : INV_X1 port map( A => registers_7_4_port, ZN => n2260);
   U2087 : INV_X1 port map( A => registers_18_5_port, ZN => n2451);
   U2088 : INV_X1 port map( A => registers_20_5_port, ZN => n2515);
   U2089 : INV_X1 port map( A => registers_26_5_port, ZN => n2579);
   U2090 : INV_X1 port map( A => registers_28_5_port, ZN => n2643);
   U2091 : INV_X1 port map( A => registers_7_5_port, ZN => n2259);
   U2092 : INV_X1 port map( A => registers_18_6_port, ZN => n2450);
   U2093 : INV_X1 port map( A => registers_20_6_port, ZN => n2514);
   U2094 : INV_X1 port map( A => registers_26_6_port, ZN => n2578);
   U2095 : INV_X1 port map( A => registers_28_6_port, ZN => n2642);
   U2096 : INV_X1 port map( A => registers_7_6_port, ZN => n2258);
   U2097 : INV_X1 port map( A => registers_18_7_port, ZN => n2449);
   U2098 : INV_X1 port map( A => registers_20_7_port, ZN => n2513);
   U2099 : INV_X1 port map( A => registers_26_7_port, ZN => n2577);
   U2100 : INV_X1 port map( A => registers_28_7_port, ZN => n2641);
   U2101 : INV_X1 port map( A => registers_7_7_port, ZN => n2257);
   U2102 : INV_X1 port map( A => registers_18_8_port, ZN => n2448);
   U2103 : INV_X1 port map( A => registers_20_8_port, ZN => n2512);
   U2104 : INV_X1 port map( A => registers_26_8_port, ZN => n2576);
   U2105 : INV_X1 port map( A => registers_28_8_port, ZN => n2640);
   U2106 : INV_X1 port map( A => registers_7_8_port, ZN => n2256);
   U2107 : INV_X1 port map( A => registers_18_9_port, ZN => n2447);
   U2108 : INV_X1 port map( A => registers_20_9_port, ZN => n2511);
   U2109 : INV_X1 port map( A => registers_26_9_port, ZN => n2575);
   U2110 : INV_X1 port map( A => registers_28_9_port, ZN => n2639);
   U2111 : INV_X1 port map( A => registers_7_9_port, ZN => n2255);
   U2112 : INV_X1 port map( A => registers_18_10_port, ZN => n2446);
   U2113 : INV_X1 port map( A => registers_20_10_port, ZN => n2510);
   U2114 : INV_X1 port map( A => registers_26_10_port, ZN => n2574);
   U2115 : INV_X1 port map( A => registers_28_10_port, ZN => n2638);
   U2116 : INV_X1 port map( A => registers_7_10_port, ZN => n2254);
   U2117 : INV_X1 port map( A => registers_18_11_port, ZN => n2445);
   U2118 : INV_X1 port map( A => registers_20_11_port, ZN => n2509);
   U2119 : INV_X1 port map( A => registers_26_11_port, ZN => n2573);
   U2120 : INV_X1 port map( A => registers_28_11_port, ZN => n2637);
   U2121 : INV_X1 port map( A => registers_7_11_port, ZN => n2253);
   U2122 : INV_X1 port map( A => registers_18_12_port, ZN => n2444);
   U2123 : INV_X1 port map( A => registers_20_12_port, ZN => n2508);
   U2124 : INV_X1 port map( A => registers_26_12_port, ZN => n2572);
   U2125 : INV_X1 port map( A => registers_28_12_port, ZN => n2636);
   U2126 : INV_X1 port map( A => registers_7_12_port, ZN => n2252);
   U2127 : INV_X1 port map( A => registers_18_13_port, ZN => n2443);
   U2128 : INV_X1 port map( A => registers_20_13_port, ZN => n2507);
   U2129 : INV_X1 port map( A => registers_26_13_port, ZN => n2571);
   U2130 : INV_X1 port map( A => registers_28_13_port, ZN => n2635);
   U2131 : INV_X1 port map( A => registers_7_13_port, ZN => n2251);
   U2132 : INV_X1 port map( A => registers_18_14_port, ZN => n2442);
   U2133 : INV_X1 port map( A => registers_20_14_port, ZN => n2506);
   U2134 : INV_X1 port map( A => registers_26_14_port, ZN => n2570);
   U2135 : INV_X1 port map( A => registers_28_14_port, ZN => n2634);
   U2136 : INV_X1 port map( A => registers_7_14_port, ZN => n2250);
   U2137 : INV_X1 port map( A => registers_18_15_port, ZN => n2441);
   U2138 : INV_X1 port map( A => registers_20_15_port, ZN => n2505);
   U2139 : INV_X1 port map( A => registers_26_15_port, ZN => n2569);
   U2140 : INV_X1 port map( A => registers_28_15_port, ZN => n2633);
   U2141 : INV_X1 port map( A => registers_7_15_port, ZN => n2249);
   U2142 : INV_X1 port map( A => registers_18_16_port, ZN => n2440);
   U2143 : INV_X1 port map( A => registers_20_16_port, ZN => n2504);
   U2144 : INV_X1 port map( A => registers_26_16_port, ZN => n2568);
   U2145 : INV_X1 port map( A => registers_28_16_port, ZN => n2632);
   U2146 : INV_X1 port map( A => registers_7_16_port, ZN => n2248);
   U2147 : INV_X1 port map( A => registers_18_17_port, ZN => n2439);
   U2148 : INV_X1 port map( A => registers_20_17_port, ZN => n2503);
   U2149 : INV_X1 port map( A => registers_26_17_port, ZN => n2567);
   U2150 : INV_X1 port map( A => registers_28_17_port, ZN => n2631);
   U2151 : INV_X1 port map( A => registers_7_17_port, ZN => n2247);
   U2152 : INV_X1 port map( A => registers_18_18_port, ZN => n2438);
   U2153 : INV_X1 port map( A => registers_20_18_port, ZN => n2502);
   U2154 : INV_X1 port map( A => registers_26_18_port, ZN => n2566);
   U2155 : INV_X1 port map( A => registers_28_18_port, ZN => n2630);
   U2156 : INV_X1 port map( A => registers_7_18_port, ZN => n2246);
   U2157 : INV_X1 port map( A => registers_18_19_port, ZN => n2437);
   U2158 : INV_X1 port map( A => registers_20_19_port, ZN => n2501);
   U2159 : INV_X1 port map( A => registers_26_19_port, ZN => n2565);
   U2160 : INV_X1 port map( A => registers_28_19_port, ZN => n2629);
   U2161 : INV_X1 port map( A => registers_7_19_port, ZN => n2245);
   U2162 : INV_X1 port map( A => registers_18_20_port, ZN => n2436);
   U2163 : INV_X1 port map( A => registers_20_20_port, ZN => n2500);
   U2164 : INV_X1 port map( A => registers_26_20_port, ZN => n2564);
   U2165 : INV_X1 port map( A => registers_28_20_port, ZN => n2628);
   U2166 : INV_X1 port map( A => registers_7_20_port, ZN => n2244);
   U2167 : INV_X1 port map( A => registers_18_21_port, ZN => n2435);
   U2168 : INV_X1 port map( A => registers_20_21_port, ZN => n2499);
   U2169 : INV_X1 port map( A => registers_26_21_port, ZN => n2563);
   U2170 : INV_X1 port map( A => registers_28_21_port, ZN => n2627);
   U2171 : INV_X1 port map( A => registers_7_21_port, ZN => n2243);
   U2172 : INV_X1 port map( A => registers_18_22_port, ZN => n2434);
   U2173 : INV_X1 port map( A => registers_20_22_port, ZN => n2498);
   U2174 : INV_X1 port map( A => registers_26_22_port, ZN => n2562);
   U2175 : INV_X1 port map( A => registers_28_22_port, ZN => n2626);
   U2176 : INV_X1 port map( A => registers_7_22_port, ZN => n2242);
   U2177 : INV_X1 port map( A => registers_18_23_port, ZN => n2433);
   U2178 : INV_X1 port map( A => registers_20_23_port, ZN => n2497);
   U2179 : INV_X1 port map( A => registers_26_23_port, ZN => n2561);
   U2180 : INV_X1 port map( A => registers_28_23_port, ZN => n2625);
   U2181 : INV_X1 port map( A => registers_7_23_port, ZN => n2241);
   U2182 : INV_X1 port map( A => registers_18_24_port, ZN => n2432);
   U2183 : INV_X1 port map( A => registers_20_24_port, ZN => n2496);
   U2184 : INV_X1 port map( A => registers_26_24_port, ZN => n2560);
   U2185 : INV_X1 port map( A => registers_28_24_port, ZN => n2624);
   U2186 : INV_X1 port map( A => registers_7_24_port, ZN => n2240);
   U2187 : INV_X1 port map( A => registers_18_25_port, ZN => n2431);
   U2188 : INV_X1 port map( A => registers_20_25_port, ZN => n2495);
   U2189 : INV_X1 port map( A => registers_26_25_port, ZN => n2559);
   U2190 : INV_X1 port map( A => registers_28_25_port, ZN => n2623);
   U2191 : INV_X1 port map( A => registers_7_25_port, ZN => n2239);
   U2192 : INV_X1 port map( A => registers_18_26_port, ZN => n2430);
   U2193 : INV_X1 port map( A => registers_20_26_port, ZN => n2494);
   U2194 : INV_X1 port map( A => registers_26_26_port, ZN => n2558);
   U2195 : INV_X1 port map( A => registers_28_26_port, ZN => n2622);
   U2196 : INV_X1 port map( A => registers_7_26_port, ZN => n2238);
   U2197 : INV_X1 port map( A => registers_18_27_port, ZN => n2429);
   U2198 : INV_X1 port map( A => registers_20_27_port, ZN => n2493);
   U2199 : INV_X1 port map( A => registers_26_27_port, ZN => n2557);
   U2200 : INV_X1 port map( A => registers_28_27_port, ZN => n2621);
   U2201 : INV_X1 port map( A => registers_7_27_port, ZN => n2237);
   U2202 : INV_X1 port map( A => registers_18_28_port, ZN => n2428);
   U2203 : INV_X1 port map( A => registers_20_28_port, ZN => n2492);
   U2204 : INV_X1 port map( A => registers_26_28_port, ZN => n2556);
   U2205 : INV_X1 port map( A => registers_28_28_port, ZN => n2620);
   U2206 : INV_X1 port map( A => registers_7_28_port, ZN => n2236);
   U2207 : INV_X1 port map( A => registers_18_29_port, ZN => n2427);
   U2208 : INV_X1 port map( A => registers_20_29_port, ZN => n2491);
   U2209 : INV_X1 port map( A => registers_26_29_port, ZN => n2555);
   U2210 : INV_X1 port map( A => registers_28_29_port, ZN => n2619);
   U2211 : INV_X1 port map( A => registers_7_29_port, ZN => n2235);
   U2212 : INV_X1 port map( A => registers_18_30_port, ZN => n2426);
   U2213 : INV_X1 port map( A => registers_20_30_port, ZN => n2490);
   U2214 : INV_X1 port map( A => registers_26_30_port, ZN => n2554);
   U2215 : INV_X1 port map( A => registers_28_30_port, ZN => n2618);
   U2216 : INV_X1 port map( A => registers_7_30_port, ZN => n2234);
   U2217 : INV_X1 port map( A => registers_18_31_port, ZN => n2425);
   U2218 : INV_X1 port map( A => registers_20_31_port, ZN => n2489);
   U2219 : INV_X1 port map( A => registers_26_31_port, ZN => n2553);
   U2220 : INV_X1 port map( A => registers_28_31_port, ZN => n2617);
   U2221 : INV_X1 port map( A => registers_7_31_port, ZN => n2233);
   U2222 : INV_X1 port map( A => add_wr(4), ZN => n2164);
   U2223 : INV_X1 port map( A => add_wr(3), ZN => n2165);
   U2224 : AND2_X1 port map( A1 => wr, A2 => n2689, ZN => n535);
   U2225 : INV_X1 port map( A => enable, ZN => n2689);
   U2226 : CLKBUF_X1 port map( A => N371, Z => n1962);
   U2227 : CLKBUF_X1 port map( A => N371, Z => n1963);
   U2228 : CLKBUF_X1 port map( A => N371, Z => n1964);
   U2229 : CLKBUF_X1 port map( A => N371, Z => n1965);
   U2230 : CLKBUF_X1 port map( A => N371, Z => n1966);
   U2231 : CLKBUF_X1 port map( A => N371, Z => n1967);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity sign_extension_sign_init26_sign_ext32 is

   port( data_in : in std_logic_vector (25 downto 0);  data_out : out 
         std_logic_vector (31 downto 0));

end sign_extension_sign_init26_sign_ext32;

architecture SYN_BEH of sign_extension_sign_init26_sign_ext32 is

begin
   data_out <= ( data_in(25), data_in(25), data_in(25), data_in(25), 
      data_in(25), data_in(25), data_in(25), data_in(24), data_in(23), 
      data_in(22), data_in(21), data_in(20), data_in(19), data_in(18), 
      data_in(17), data_in(16), data_in(15), data_in(14), data_in(13), 
      data_in(12), data_in(11), data_in(10), data_in(9), data_in(8), data_in(7)
      , data_in(6), data_in(5), data_in(4), data_in(3), data_in(2), data_in(1),
      data_in(0) );

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_17 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_17;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_17 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42
      , n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n49, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n49, Q => Q(30), 
                           QN => n67);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n49, Q => Q(29), 
                           QN => n68);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n49, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n49, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n49, Q => Q(26), 
                           QN => n71);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n49, Q => Q(25), 
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n49, Q => Q(24), 
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n48, Q => Q(23), 
                           QN => n74);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n48, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n48, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n48, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n48, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n48, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n48, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n48, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n48, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n48, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n48, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n48, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n47, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n47, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n47, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n47, Q => Q(8), 
                           QN => n89);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n47, Q => Q(7), 
                           QN => n90);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n47, Q => Q(6), 
                           QN => n91);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n47, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n47, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n47, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n47, Q => Q(2), 
                           QN => n95);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n47, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n47, Q => Q(0), 
                           QN => n97);
   U2 : BUF_X1 port map( A => RESET_n, Z => n47);
   U3 : BUF_X1 port map( A => RESET_n, Z => n48);
   U4 : BUF_X1 port map( A => RESET_n, Z => n49);
   U5 : INV_X1 port map( A => n46, ZN => n37);
   U6 : INV_X1 port map( A => n46, ZN => n36);
   U7 : BUF_X1 port map( A => n35, Z => n46);
   U8 : BUF_X1 port map( A => n34, Z => n41);
   U9 : BUF_X1 port map( A => n34, Z => n42);
   U10 : BUF_X1 port map( A => n35, Z => n44);
   U11 : BUF_X1 port map( A => n33, Z => n38);
   U12 : BUF_X1 port map( A => n33, Z => n39);
   U13 : BUF_X1 port map( A => n33, Z => n40);
   U14 : BUF_X1 port map( A => n34, Z => n43);
   U15 : BUF_X1 port map( A => n35, Z => n45);
   U16 : OAI22_X1 port map( A1 => n97, A2 => n37, B1 => n39, B2 => n113, ZN => 
                           n32);
   U17 : INV_X1 port map( A => D(0), ZN => n113);
   U18 : OAI22_X1 port map( A1 => n96, A2 => n36, B1 => n39, B2 => n112, ZN => 
                           n31);
   U19 : INV_X1 port map( A => D(1), ZN => n112);
   U20 : OAI22_X1 port map( A1 => n95, A2 => n37, B1 => n40, B2 => n111, ZN => 
                           n30);
   U21 : INV_X1 port map( A => D(2), ZN => n111);
   U22 : OAI22_X1 port map( A1 => n94, A2 => n37, B1 => n40, B2 => n110, ZN => 
                           n29);
   U23 : INV_X1 port map( A => D(3), ZN => n110);
   U24 : OAI22_X1 port map( A1 => n93, A2 => n37, B1 => n40, B2 => n109, ZN => 
                           n28);
   U25 : INV_X1 port map( A => D(4), ZN => n109);
   U26 : OAI22_X1 port map( A1 => n92, A2 => n37, B1 => n41, B2 => n108, ZN => 
                           n27);
   U27 : INV_X1 port map( A => D(5), ZN => n108);
   U28 : OAI22_X1 port map( A1 => n91, A2 => n37, B1 => n41, B2 => n107, ZN => 
                           n26);
   U29 : INV_X1 port map( A => D(6), ZN => n107);
   U30 : OAI22_X1 port map( A1 => n90, A2 => n37, B1 => n41, B2 => n106, ZN => 
                           n25);
   U31 : INV_X1 port map( A => D(7), ZN => n106);
   U32 : OAI22_X1 port map( A1 => n89, A2 => n37, B1 => n41, B2 => n105, ZN => 
                           n24);
   U33 : INV_X1 port map( A => D(8), ZN => n105);
   U34 : OAI22_X1 port map( A1 => n88, A2 => n37, B1 => n42, B2 => n104, ZN => 
                           n23);
   U35 : INV_X1 port map( A => D(9), ZN => n104);
   U36 : OAI22_X1 port map( A1 => n87, A2 => n37, B1 => n42, B2 => n103, ZN => 
                           n22);
   U37 : INV_X1 port map( A => D(10), ZN => n103);
   U38 : OAI22_X1 port map( A1 => n86, A2 => n37, B1 => n42, B2 => n102, ZN => 
                           n21);
   U39 : INV_X1 port map( A => D(11), ZN => n102);
   U40 : OAI22_X1 port map( A1 => n85, A2 => n37, B1 => n42, B2 => n101, ZN => 
                           n20);
   U41 : INV_X1 port map( A => D(12), ZN => n101);
   U42 : OAI22_X1 port map( A1 => n84, A2 => n36, B1 => n43, B2 => n100, ZN => 
                           n19);
   U43 : INV_X1 port map( A => D(13), ZN => n100);
   U44 : OAI22_X1 port map( A1 => n83, A2 => n36, B1 => n43, B2 => n99, ZN => 
                           n18);
   U45 : INV_X1 port map( A => D(14), ZN => n99);
   U46 : OAI22_X1 port map( A1 => n82, A2 => n36, B1 => n43, B2 => n98, ZN => 
                           n17);
   U47 : INV_X1 port map( A => D(15), ZN => n98);
   U48 : OAI22_X1 port map( A1 => n81, A2 => n36, B1 => n44, B2 => n65, ZN => 
                           n16);
   U49 : INV_X1 port map( A => D(16), ZN => n65);
   U50 : OAI22_X1 port map( A1 => n80, A2 => n36, B1 => n44, B2 => n64, ZN => 
                           n15);
   U51 : INV_X1 port map( A => D(17), ZN => n64);
   U52 : OAI22_X1 port map( A1 => n79, A2 => n36, B1 => n44, B2 => n63, ZN => 
                           n14);
   U53 : INV_X1 port map( A => D(18), ZN => n63);
   U54 : OAI22_X1 port map( A1 => n78, A2 => n36, B1 => n44, B2 => n62, ZN => 
                           n13);
   U55 : INV_X1 port map( A => D(19), ZN => n62);
   U56 : OAI22_X1 port map( A1 => n77, A2 => n36, B1 => n45, B2 => n61, ZN => 
                           n12);
   U57 : INV_X1 port map( A => D(20), ZN => n61);
   U58 : OAI22_X1 port map( A1 => n76, A2 => n36, B1 => n45, B2 => n60, ZN => 
                           n11);
   U59 : INV_X1 port map( A => D(21), ZN => n60);
   U60 : OAI22_X1 port map( A1 => n75, A2 => n36, B1 => n45, B2 => n59, ZN => 
                           n10);
   U61 : INV_X1 port map( A => D(22), ZN => n59);
   U62 : OAI22_X1 port map( A1 => n74, A2 => n37, B1 => n38, B2 => n58, ZN => 
                           n9);
   U63 : INV_X1 port map( A => D(23), ZN => n58);
   U64 : OAI22_X1 port map( A1 => n73, A2 => n36, B1 => n38, B2 => n57, ZN => 
                           n8);
   U65 : INV_X1 port map( A => D(24), ZN => n57);
   U66 : OAI22_X1 port map( A1 => n72, A2 => n37, B1 => n38, B2 => n56, ZN => 
                           n7);
   U67 : INV_X1 port map( A => D(25), ZN => n56);
   U68 : OAI22_X1 port map( A1 => n71, A2 => n36, B1 => n38, B2 => n55, ZN => 
                           n6);
   U69 : INV_X1 port map( A => D(26), ZN => n55);
   U70 : OAI22_X1 port map( A1 => n70, A2 => n37, B1 => n39, B2 => n54, ZN => 
                           n5);
   U71 : INV_X1 port map( A => D(27), ZN => n54);
   U72 : OAI22_X1 port map( A1 => n69, A2 => n36, B1 => n39, B2 => n53, ZN => 
                           n4);
   U73 : INV_X1 port map( A => D(28), ZN => n53);
   U74 : OAI22_X1 port map( A1 => n68, A2 => n37, B1 => n40, B2 => n52, ZN => 
                           n3);
   U75 : INV_X1 port map( A => D(29), ZN => n52);
   U76 : OAI22_X1 port map( A1 => n67, A2 => n36, B1 => n43, B2 => n51, ZN => 
                           n2);
   U77 : INV_X1 port map( A => D(30), ZN => n51);
   U78 : OAI22_X1 port map( A1 => n66, A2 => n36, B1 => n45, B2 => n50, ZN => 
                           n1);
   U79 : INV_X1 port map( A => D(31), ZN => n50);
   U80 : BUF_X1 port map( A => Enable_n, Z => n35);
   U81 : BUF_X1 port map( A => Enable_n, Z => n33);
   U82 : BUF_X1 port map( A => Enable_n, Z => n34);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_18 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_18;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_18 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n47, Q => Q(31), 
                           QN => n145);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n47, Q => Q(30), 
                           QN => n144);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n47, Q => Q(29), 
                           QN => n143);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n47, Q => Q(28), 
                           QN => n142);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n47, Q => Q(27), 
                           QN => n141);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n47, Q => Q(26), 
                           QN => n140);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n47, Q => Q(25), 
                           QN => n139);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n47, Q => Q(24), 
                           QN => n138);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n47, Q => Q(23), 
                           QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n47, Q => Q(22),
                           QN => n136);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n47, Q => Q(21),
                           QN => n135);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n47, Q => Q(20),
                           QN => n134);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n48, Q => Q(19),
                           QN => n133);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n48, Q => Q(18),
                           QN => n132);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n48, Q => Q(17),
                           QN => n131);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n48, Q => Q(16),
                           QN => n130);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n48, Q => Q(15),
                           QN => n129);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n48, Q => Q(14),
                           QN => n128);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n48, Q => Q(13),
                           QN => n127);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n48, Q => Q(12),
                           QN => n126);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n48, Q => Q(11),
                           QN => n125);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n48, Q => Q(10),
                           QN => n124);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n48, Q => Q(9), 
                           QN => n123);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n48, Q => Q(8), 
                           QN => n122);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n49, Q => Q(7), 
                           QN => n121);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n49, Q => Q(6), 
                           QN => n120);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n49, Q => Q(5), 
                           QN => n119);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n49, Q => Q(4), 
                           QN => n118);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n49, Q => Q(3), 
                           QN => n117);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n49, Q => Q(2), 
                           QN => n116);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n49, Q => Q(1), 
                           QN => n115);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n49, Q => Q(0), 
                           QN => n114);
   U2 : BUF_X1 port map( A => RESET_n, Z => n48);
   U3 : BUF_X1 port map( A => RESET_n, Z => n47);
   U4 : BUF_X1 port map( A => RESET_n, Z => n49);
   U5 : INV_X1 port map( A => n46, ZN => n37);
   U6 : INV_X1 port map( A => n46, ZN => n36);
   U7 : BUF_X1 port map( A => n35, Z => n46);
   U8 : BUF_X1 port map( A => n34, Z => n41);
   U9 : BUF_X1 port map( A => n34, Z => n42);
   U10 : BUF_X1 port map( A => n35, Z => n44);
   U11 : BUF_X1 port map( A => n33, Z => n38);
   U12 : BUF_X1 port map( A => n33, Z => n39);
   U13 : BUF_X1 port map( A => n33, Z => n40);
   U14 : BUF_X1 port map( A => n34, Z => n43);
   U15 : BUF_X1 port map( A => n35, Z => n45);
   U16 : OAI22_X1 port map( A1 => n114, A2 => n37, B1 => n39, B2 => n113, ZN =>
                           n32);
   U17 : INV_X1 port map( A => D(0), ZN => n113);
   U18 : OAI22_X1 port map( A1 => n115, A2 => n36, B1 => n39, B2 => n112, ZN =>
                           n31);
   U19 : INV_X1 port map( A => D(1), ZN => n112);
   U20 : OAI22_X1 port map( A1 => n116, A2 => n37, B1 => n40, B2 => n111, ZN =>
                           n30);
   U21 : INV_X1 port map( A => D(2), ZN => n111);
   U22 : OAI22_X1 port map( A1 => n117, A2 => n37, B1 => n40, B2 => n110, ZN =>
                           n29);
   U23 : INV_X1 port map( A => D(3), ZN => n110);
   U24 : OAI22_X1 port map( A1 => n134, A2 => n36, B1 => n45, B2 => n65, ZN => 
                           n12);
   U25 : INV_X1 port map( A => D(20), ZN => n65);
   U26 : OAI22_X1 port map( A1 => n135, A2 => n36, B1 => n45, B2 => n64, ZN => 
                           n11);
   U27 : INV_X1 port map( A => D(21), ZN => n64);
   U28 : OAI22_X1 port map( A1 => n136, A2 => n36, B1 => n45, B2 => n63, ZN => 
                           n10);
   U29 : INV_X1 port map( A => D(22), ZN => n63);
   U30 : OAI22_X1 port map( A1 => n137, A2 => n37, B1 => n38, B2 => n62, ZN => 
                           n9);
   U31 : INV_X1 port map( A => D(23), ZN => n62);
   U32 : OAI22_X1 port map( A1 => n138, A2 => n37, B1 => n38, B2 => n101, ZN =>
                           n8);
   U33 : INV_X1 port map( A => D(24), ZN => n101);
   U34 : OAI22_X1 port map( A1 => n139, A2 => n36, B1 => n38, B2 => n100, ZN =>
                           n7);
   U35 : INV_X1 port map( A => D(25), ZN => n100);
   U36 : OAI22_X1 port map( A1 => n140, A2 => n37, B1 => n38, B2 => n99, ZN => 
                           n6);
   U37 : INV_X1 port map( A => D(26), ZN => n99);
   U38 : OAI22_X1 port map( A1 => n141, A2 => n36, B1 => n39, B2 => n98, ZN => 
                           n5);
   U39 : INV_X1 port map( A => D(27), ZN => n98);
   U40 : OAI22_X1 port map( A1 => n142, A2 => n36, B1 => n39, B2 => n105, ZN =>
                           n4);
   U41 : INV_X1 port map( A => D(28), ZN => n105);
   U42 : OAI22_X1 port map( A1 => n143, A2 => n37, B1 => n40, B2 => n104, ZN =>
                           n3);
   U43 : INV_X1 port map( A => D(29), ZN => n104);
   U44 : OAI22_X1 port map( A1 => n144, A2 => n36, B1 => n43, B2 => n103, ZN =>
                           n2);
   U45 : INV_X1 port map( A => D(30), ZN => n103);
   U46 : OAI22_X1 port map( A1 => n145, A2 => n36, B1 => n45, B2 => n102, ZN =>
                           n1);
   U47 : INV_X1 port map( A => D(31), ZN => n102);
   U48 : OAI22_X1 port map( A1 => n130, A2 => n36, B1 => n44, B2 => n61, ZN => 
                           n16);
   U49 : INV_X1 port map( A => D(16), ZN => n61);
   U50 : OAI22_X1 port map( A1 => n131, A2 => n36, B1 => n44, B2 => n60, ZN => 
                           n15);
   U51 : INV_X1 port map( A => D(17), ZN => n60);
   U52 : OAI22_X1 port map( A1 => n132, A2 => n36, B1 => n44, B2 => n59, ZN => 
                           n14);
   U53 : INV_X1 port map( A => D(18), ZN => n59);
   U54 : OAI22_X1 port map( A1 => n122, A2 => n37, B1 => n41, B2 => n53, ZN => 
                           n24);
   U55 : INV_X1 port map( A => D(8), ZN => n53);
   U56 : OAI22_X1 port map( A1 => n123, A2 => n37, B1 => n42, B2 => n52, ZN => 
                           n23);
   U57 : INV_X1 port map( A => D(9), ZN => n52);
   U58 : OAI22_X1 port map( A1 => n124, A2 => n37, B1 => n42, B2 => n51, ZN => 
                           n22);
   U59 : INV_X1 port map( A => D(10), ZN => n51);
   U60 : OAI22_X1 port map( A1 => n133, A2 => n36, B1 => n44, B2 => n58, ZN => 
                           n13);
   U61 : INV_X1 port map( A => D(19), ZN => n58);
   U62 : OAI22_X1 port map( A1 => n118, A2 => n37, B1 => n40, B2 => n109, ZN =>
                           n28);
   U63 : INV_X1 port map( A => D(4), ZN => n109);
   U64 : OAI22_X1 port map( A1 => n119, A2 => n37, B1 => n41, B2 => n108, ZN =>
                           n27);
   U65 : INV_X1 port map( A => D(5), ZN => n108);
   U66 : OAI22_X1 port map( A1 => n120, A2 => n37, B1 => n41, B2 => n107, ZN =>
                           n26);
   U67 : INV_X1 port map( A => D(6), ZN => n107);
   U68 : OAI22_X1 port map( A1 => n126, A2 => n37, B1 => n42, B2 => n57, ZN => 
                           n20);
   U69 : INV_X1 port map( A => D(12), ZN => n57);
   U70 : OAI22_X1 port map( A1 => n127, A2 => n36, B1 => n43, B2 => n56, ZN => 
                           n19);
   U71 : INV_X1 port map( A => D(13), ZN => n56);
   U72 : OAI22_X1 port map( A1 => n128, A2 => n36, B1 => n43, B2 => n55, ZN => 
                           n18);
   U73 : INV_X1 port map( A => D(14), ZN => n55);
   U74 : OAI22_X1 port map( A1 => n125, A2 => n37, B1 => n42, B2 => n50, ZN => 
                           n21);
   U75 : INV_X1 port map( A => D(11), ZN => n50);
   U76 : OAI22_X1 port map( A1 => n121, A2 => n37, B1 => n41, B2 => n106, ZN =>
                           n25);
   U77 : INV_X1 port map( A => D(7), ZN => n106);
   U78 : OAI22_X1 port map( A1 => n129, A2 => n36, B1 => n43, B2 => n54, ZN => 
                           n17);
   U79 : INV_X1 port map( A => D(15), ZN => n54);
   U80 : BUF_X1 port map( A => Enable_n, Z => n35);
   U81 : BUF_X1 port map( A => Enable_n, Z => n33);
   U82 : BUF_X1 port map( A => Enable_n, Z => n34);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity P4_ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic;  Y : out std_logic_vector (31 downto 0));

end P4_ADDER_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32_NBIT_PER_BLOCK4_0 is

   component SUMGEN_NBIT32_NBLOCKS8_0
      port( A, B : in std_logic_vector (31 downto 0);  cin_vect : in 
            std_logic_vector (7 downto 0);  Co : out std_logic;  SUM : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal outCarryGen_7_port, outCarryGen_6_port, outCarryGen_5_port, 
      outCarryGen_4_port, outCarryGen_3_port, outCarryGen_2_port, 
      outCarryGen_1_port, outCarryGen_0_port : std_logic;

begin
   
   CG : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Cin => Cin, Co(7) 
                           => outCarryGen_7_port, Co(6) => outCarryGen_6_port, 
                           Co(5) => outCarryGen_5_port, Co(4) => 
                           outCarryGen_4_port, Co(3) => outCarryGen_3_port, 
                           Co(2) => outCarryGen_2_port, Co(1) => 
                           outCarryGen_1_port, Co(0) => outCarryGen_0_port);
   SG : SUMGEN_NBIT32_NBLOCKS8_0 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), cin_vect(7) => 
                           outCarryGen_7_port, cin_vect(6) => 
                           outCarryGen_6_port, cin_vect(5) => 
                           outCarryGen_5_port, cin_vect(4) => 
                           outCarryGen_4_port, cin_vect(3) => 
                           outCarryGen_3_port, cin_vect(2) => 
                           outCarryGen_2_port, cin_vect(1) => 
                           outCarryGen_1_port, cin_vect(0) => 
                           outCarryGen_0_port, Co => Cout, SUM(31) => Y(31), 
                           SUM(30) => Y(30), SUM(29) => Y(29), SUM(28) => Y(28)
                           , SUM(27) => Y(27), SUM(26) => Y(26), SUM(25) => 
                           Y(25), SUM(24) => Y(24), SUM(23) => Y(23), SUM(22) 
                           => Y(22), SUM(21) => Y(21), SUM(20) => Y(20), 
                           SUM(19) => Y(19), SUM(18) => Y(18), SUM(17) => Y(17)
                           , SUM(16) => Y(16), SUM(15) => Y(15), SUM(14) => 
                           Y(14), SUM(13) => Y(13), SUM(12) => Y(12), SUM(11) 
                           => Y(11), SUM(10) => Y(10), SUM(9) => Y(9), SUM(8) 
                           => Y(8), SUM(7) => Y(7), SUM(6) => Y(6), SUM(5) => 
                           Y(5), SUM(4) => Y(4), SUM(3) => Y(3), SUM(2) => Y(2)
                           , SUM(1) => Y(1), SUM(0) => Y(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity REG_GEN_NBIT32_0 is

   port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end REG_GEN_NBIT32_0;

architecture SYN_REG_ASYNCH of REG_GEN_NBIT32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42
      , n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n47, Q => Q(31), 
                           QN => n66);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n47, Q => Q(30), 
                           QN => n67);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n47, Q => Q(29), 
                           QN => n68);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n47, Q => Q(28), 
                           QN => n69);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n47, Q => Q(27), 
                           QN => n70);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n47, Q => Q(26), 
                           QN => n71);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n47, Q => Q(25), 
                           QN => n72);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n47, Q => Q(24), 
                           QN => n73);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n47, Q => Q(23), 
                           QN => n74);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n47, Q => Q(22),
                           QN => n75);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n47, Q => Q(21),
                           QN => n76);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n47, Q => Q(20),
                           QN => n77);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n48, Q => Q(19),
                           QN => n78);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n48, Q => Q(18),
                           QN => n79);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n48, Q => Q(17),
                           QN => n80);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n48, Q => Q(16),
                           QN => n81);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n48, Q => Q(15),
                           QN => n82);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n48, Q => Q(14),
                           QN => n83);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n48, Q => Q(13),
                           QN => n84);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n48, Q => Q(12),
                           QN => n85);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n48, Q => Q(11),
                           QN => n86);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n48, Q => Q(10),
                           QN => n87);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n48, Q => Q(9), 
                           QN => n88);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n48, Q => Q(8), 
                           QN => n89);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n49, Q => Q(7), 
                           QN => n90);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n49, Q => Q(6), 
                           QN => n91);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n49, Q => Q(5), 
                           QN => n92);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n49, Q => Q(4), 
                           QN => n93);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n49, Q => Q(3), 
                           QN => n94);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n49, Q => Q(2), 
                           QN => n95);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n49, Q => Q(1), 
                           QN => n96);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n49, Q => Q(0), 
                           QN => n97);
   U2 : BUF_X1 port map( A => RESET_n, Z => n48);
   U3 : BUF_X1 port map( A => RESET_n, Z => n47);
   U4 : BUF_X1 port map( A => RESET_n, Z => n49);
   U5 : INV_X1 port map( A => n46, ZN => n37);
   U6 : INV_X1 port map( A => n46, ZN => n36);
   U7 : BUF_X1 port map( A => n35, Z => n46);
   U8 : BUF_X1 port map( A => n34, Z => n41);
   U9 : BUF_X1 port map( A => n34, Z => n42);
   U10 : BUF_X1 port map( A => n35, Z => n44);
   U11 : BUF_X1 port map( A => n33, Z => n38);
   U12 : BUF_X1 port map( A => n33, Z => n39);
   U13 : BUF_X1 port map( A => n33, Z => n40);
   U14 : BUF_X1 port map( A => n34, Z => n43);
   U15 : BUF_X1 port map( A => n35, Z => n45);
   U16 : OAI22_X1 port map( A1 => n85, A2 => n37, B1 => n42, B2 => n57, ZN => 
                           n20);
   U17 : INV_X1 port map( A => D(12), ZN => n57);
   U18 : OAI22_X1 port map( A1 => n84, A2 => n36, B1 => n43, B2 => n56, ZN => 
                           n19);
   U19 : INV_X1 port map( A => D(13), ZN => n56);
   U20 : OAI22_X1 port map( A1 => n82, A2 => n36, B1 => n43, B2 => n54, ZN => 
                           n17);
   U21 : INV_X1 port map( A => D(15), ZN => n54);
   U22 : OAI22_X1 port map( A1 => n81, A2 => n36, B1 => n44, B2 => n61, ZN => 
                           n16);
   U23 : INV_X1 port map( A => D(16), ZN => n61);
   U24 : OAI22_X1 port map( A1 => n79, A2 => n36, B1 => n44, B2 => n59, ZN => 
                           n14);
   U25 : INV_X1 port map( A => D(18), ZN => n59);
   U26 : OAI22_X1 port map( A1 => n78, A2 => n36, B1 => n44, B2 => n58, ZN => 
                           n13);
   U27 : INV_X1 port map( A => D(19), ZN => n58);
   U28 : OAI22_X1 port map( A1 => n77, A2 => n36, B1 => n45, B2 => n65, ZN => 
                           n12);
   U29 : INV_X1 port map( A => D(20), ZN => n65);
   U30 : OAI22_X1 port map( A1 => n75, A2 => n36, B1 => n45, B2 => n63, ZN => 
                           n10);
   U31 : INV_X1 port map( A => D(22), ZN => n63);
   U32 : OAI22_X1 port map( A1 => n74, A2 => n37, B1 => n38, B2 => n62, ZN => 
                           n9);
   U33 : INV_X1 port map( A => D(23), ZN => n62);
   U34 : OAI22_X1 port map( A1 => n73, A2 => n36, B1 => n38, B2 => n101, ZN => 
                           n8);
   U35 : INV_X1 port map( A => D(24), ZN => n101);
   U36 : OAI22_X1 port map( A1 => n72, A2 => n37, B1 => n38, B2 => n100, ZN => 
                           n7);
   U37 : INV_X1 port map( A => D(25), ZN => n100);
   U38 : OAI22_X1 port map( A1 => n71, A2 => n36, B1 => n38, B2 => n99, ZN => 
                           n6);
   U39 : INV_X1 port map( A => D(26), ZN => n99);
   U40 : OAI22_X1 port map( A1 => n70, A2 => n37, B1 => n39, B2 => n98, ZN => 
                           n5);
   U41 : INV_X1 port map( A => D(27), ZN => n98);
   U42 : OAI22_X1 port map( A1 => n69, A2 => n36, B1 => n39, B2 => n105, ZN => 
                           n4);
   U43 : INV_X1 port map( A => D(28), ZN => n105);
   U44 : OAI22_X1 port map( A1 => n68, A2 => n37, B1 => n40, B2 => n104, ZN => 
                           n3);
   U45 : INV_X1 port map( A => D(29), ZN => n104);
   U46 : OAI22_X1 port map( A1 => n67, A2 => n36, B1 => n43, B2 => n103, ZN => 
                           n2);
   U47 : INV_X1 port map( A => D(30), ZN => n103);
   U48 : OAI22_X1 port map( A1 => n66, A2 => n36, B1 => n45, B2 => n102, ZN => 
                           n1);
   U49 : INV_X1 port map( A => D(31), ZN => n102);
   U50 : OAI22_X1 port map( A1 => n83, A2 => n36, B1 => n43, B2 => n55, ZN => 
                           n18);
   U51 : INV_X1 port map( A => D(14), ZN => n55);
   U52 : OAI22_X1 port map( A1 => n80, A2 => n36, B1 => n44, B2 => n60, ZN => 
                           n15);
   U53 : INV_X1 port map( A => D(17), ZN => n60);
   U54 : OAI22_X1 port map( A1 => n76, A2 => n36, B1 => n45, B2 => n64, ZN => 
                           n11);
   U55 : INV_X1 port map( A => D(21), ZN => n64);
   U56 : OAI22_X1 port map( A1 => n90, A2 => n37, B1 => n41, B2 => n106, ZN => 
                           n25);
   U57 : INV_X1 port map( A => D(7), ZN => n106);
   U58 : OAI22_X1 port map( A1 => n94, A2 => n37, B1 => n40, B2 => n110, ZN => 
                           n29);
   U59 : INV_X1 port map( A => D(3), ZN => n110);
   U60 : OAI22_X1 port map( A1 => n97, A2 => n37, B1 => n39, B2 => n113, ZN => 
                           n32);
   U61 : INV_X1 port map( A => D(0), ZN => n113);
   U62 : OAI22_X1 port map( A1 => n96, A2 => n36, B1 => n39, B2 => n112, ZN => 
                           n31);
   U63 : INV_X1 port map( A => D(1), ZN => n112);
   U64 : OAI22_X1 port map( A1 => n95, A2 => n37, B1 => n40, B2 => n111, ZN => 
                           n30);
   U65 : INV_X1 port map( A => D(2), ZN => n111);
   U66 : OAI22_X1 port map( A1 => n93, A2 => n37, B1 => n40, B2 => n109, ZN => 
                           n28);
   U67 : INV_X1 port map( A => D(4), ZN => n109);
   U68 : OAI22_X1 port map( A1 => n92, A2 => n37, B1 => n41, B2 => n108, ZN => 
                           n27);
   U69 : INV_X1 port map( A => D(5), ZN => n108);
   U70 : OAI22_X1 port map( A1 => n91, A2 => n37, B1 => n41, B2 => n107, ZN => 
                           n26);
   U71 : INV_X1 port map( A => D(6), ZN => n107);
   U72 : OAI22_X1 port map( A1 => n89, A2 => n37, B1 => n41, B2 => n53, ZN => 
                           n24);
   U73 : INV_X1 port map( A => D(8), ZN => n53);
   U74 : OAI22_X1 port map( A1 => n87, A2 => n37, B1 => n42, B2 => n51, ZN => 
                           n22);
   U75 : INV_X1 port map( A => D(10), ZN => n51);
   U76 : OAI22_X1 port map( A1 => n86, A2 => n37, B1 => n42, B2 => n50, ZN => 
                           n21);
   U77 : INV_X1 port map( A => D(11), ZN => n50);
   U78 : OAI22_X1 port map( A1 => n88, A2 => n37, B1 => n42, B2 => n52, ZN => 
                           n23);
   U79 : INV_X1 port map( A => D(9), ZN => n52);
   U80 : BUF_X1 port map( A => Enable_n, Z => n35);
   U81 : BUF_X1 port map( A => Enable_n, Z => n33);
   U82 : BUF_X1 port map( A => Enable_n, Z => n34);

end SYN_REG_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_NBIT32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n33, n66, n67, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n100, Z => n33);
   U2 : BUF_X1 port map( A => n100, Z => n66);
   U3 : BUF_X1 port map( A => n100, Z => n67);
   U4 : INV_X1 port map( A => n62, ZN => Y(12));
   U5 : AOI22_X1 port map( A1 => A(12), A2 => n33, B1 => B(12), B2 => SEL, ZN 
                           => n62);
   U6 : INV_X1 port map( A => n61, ZN => Y(13));
   U7 : AOI22_X1 port map( A1 => A(13), A2 => n33, B1 => B(13), B2 => SEL, ZN 
                           => n61);
   U8 : INV_X1 port map( A => n59, ZN => Y(15));
   U9 : AOI22_X1 port map( A1 => A(15), A2 => n33, B1 => B(15), B2 => SEL, ZN 
                           => n59);
   U10 : INV_X1 port map( A => n58, ZN => Y(16));
   U11 : AOI22_X1 port map( A1 => A(16), A2 => n33, B1 => B(16), B2 => SEL, ZN 
                           => n58);
   U12 : INV_X1 port map( A => n56, ZN => Y(18));
   U13 : AOI22_X1 port map( A1 => A(18), A2 => n33, B1 => B(18), B2 => SEL, ZN 
                           => n56);
   U14 : INV_X1 port map( A => n55, ZN => Y(19));
   U15 : AOI22_X1 port map( A1 => A(19), A2 => n33, B1 => B(19), B2 => SEL, ZN 
                           => n55);
   U16 : INV_X1 port map( A => n53, ZN => Y(20));
   U17 : AOI22_X1 port map( A1 => A(20), A2 => n66, B1 => B(20), B2 => SEL, ZN 
                           => n53);
   U18 : INV_X1 port map( A => n51, ZN => Y(22));
   U19 : AOI22_X1 port map( A1 => A(22), A2 => n66, B1 => B(22), B2 => SEL, ZN 
                           => n51);
   U20 : INV_X1 port map( A => n50, ZN => Y(23));
   U21 : AOI22_X1 port map( A1 => A(23), A2 => n66, B1 => B(23), B2 => SEL, ZN 
                           => n50);
   U22 : INV_X1 port map( A => n49, ZN => Y(24));
   U23 : AOI22_X1 port map( A1 => A(24), A2 => n66, B1 => B(24), B2 => SEL, ZN 
                           => n49);
   U24 : INV_X1 port map( A => n48, ZN => Y(25));
   U25 : AOI22_X1 port map( A1 => A(25), A2 => n66, B1 => B(25), B2 => SEL, ZN 
                           => n48);
   U26 : INV_X1 port map( A => n47, ZN => Y(26));
   U27 : AOI22_X1 port map( A1 => A(26), A2 => n66, B1 => B(26), B2 => SEL, ZN 
                           => n47);
   U28 : INV_X1 port map( A => n46, ZN => Y(27));
   U29 : AOI22_X1 port map( A1 => A(27), A2 => n66, B1 => B(27), B2 => SEL, ZN 
                           => n46);
   U30 : INV_X1 port map( A => n45, ZN => Y(28));
   U31 : AOI22_X1 port map( A1 => A(28), A2 => n66, B1 => B(28), B2 => SEL, ZN 
                           => n45);
   U32 : INV_X1 port map( A => n44, ZN => Y(29));
   U33 : AOI22_X1 port map( A1 => A(29), A2 => n66, B1 => B(29), B2 => SEL, ZN 
                           => n44);
   U34 : INV_X1 port map( A => n42, ZN => Y(30));
   U35 : AOI22_X1 port map( A1 => A(30), A2 => n66, B1 => B(30), B2 => SEL, ZN 
                           => n42);
   U36 : INV_X1 port map( A => n41, ZN => Y(31));
   U37 : AOI22_X1 port map( A1 => A(31), A2 => n67, B1 => B(31), B2 => SEL, ZN 
                           => n41);
   U38 : INV_X1 port map( A => n60, ZN => Y(14));
   U39 : AOI22_X1 port map( A1 => A(14), A2 => n33, B1 => B(14), B2 => SEL, ZN 
                           => n60);
   U40 : INV_X1 port map( A => n57, ZN => Y(17));
   U41 : AOI22_X1 port map( A1 => A(17), A2 => n33, B1 => B(17), B2 => SEL, ZN 
                           => n57);
   U42 : INV_X1 port map( A => n52, ZN => Y(21));
   U43 : AOI22_X1 port map( A1 => A(21), A2 => n66, B1 => B(21), B2 => SEL, ZN 
                           => n52);
   U44 : INV_X1 port map( A => n36, ZN => Y(7));
   U45 : AOI22_X1 port map( A1 => A(7), A2 => n67, B1 => B(7), B2 => SEL, ZN =>
                           n36);
   U46 : INV_X1 port map( A => n40, ZN => Y(3));
   U47 : AOI22_X1 port map( A1 => A(3), A2 => n67, B1 => B(3), B2 => SEL, ZN =>
                           n40);
   U48 : INV_X1 port map( A => n65, ZN => Y(0));
   U49 : AOI22_X1 port map( A1 => A(0), A2 => n33, B1 => B(0), B2 => SEL, ZN =>
                           n65);
   U50 : INV_X1 port map( A => n54, ZN => Y(1));
   U51 : AOI22_X1 port map( A1 => A(1), A2 => n33, B1 => B(1), B2 => SEL, ZN =>
                           n54);
   U52 : INV_X1 port map( A => n43, ZN => Y(2));
   U53 : AOI22_X1 port map( A1 => A(2), A2 => n66, B1 => B(2), B2 => SEL, ZN =>
                           n43);
   U54 : INV_X1 port map( A => n39, ZN => Y(4));
   U55 : AOI22_X1 port map( A1 => A(4), A2 => n67, B1 => B(4), B2 => SEL, ZN =>
                           n39);
   U56 : INV_X1 port map( A => n38, ZN => Y(5));
   U57 : AOI22_X1 port map( A1 => A(5), A2 => n67, B1 => B(5), B2 => SEL, ZN =>
                           n38);
   U58 : INV_X1 port map( A => n37, ZN => Y(6));
   U59 : AOI22_X1 port map( A1 => A(6), A2 => n67, B1 => B(6), B2 => SEL, ZN =>
                           n37);
   U60 : INV_X1 port map( A => n35, ZN => Y(8));
   U61 : AOI22_X1 port map( A1 => A(8), A2 => n67, B1 => B(8), B2 => SEL, ZN =>
                           n35);
   U62 : INV_X1 port map( A => n64, ZN => Y(10));
   U63 : AOI22_X1 port map( A1 => A(10), A2 => n33, B1 => B(10), B2 => SEL, ZN 
                           => n64);
   U64 : INV_X1 port map( A => n63, ZN => Y(11));
   U65 : AOI22_X1 port map( A1 => A(11), A2 => n33, B1 => B(11), B2 => SEL, ZN 
                           => n63);
   U66 : INV_X1 port map( A => n34, ZN => Y(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n67, B1 => SEL, B2 => B(9), ZN =>
                           n34);
   U68 : INV_X1 port map( A => SEL, ZN => n100);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity writeBackUnit_nbit32 is

   port( MemtoReg : in std_logic;  ReadData, AluResult : in std_logic_vector 
         (31 downto 0);  WriteData : out std_logic_vector (31 downto 0));

end writeBackUnit_nbit32;

architecture SYN_struct of writeBackUnit_nbit32 is

   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;

begin
   
   mux_writeBack : MUX21_GENERIC_NBIT32_3 port map( A(31) => ReadData(31), 
                           A(30) => ReadData(30), A(29) => ReadData(29), A(28) 
                           => ReadData(28), A(27) => ReadData(27), A(26) => 
                           ReadData(26), A(25) => ReadData(25), A(24) => 
                           ReadData(24), A(23) => ReadData(23), A(22) => 
                           ReadData(22), A(21) => ReadData(21), A(20) => 
                           ReadData(20), A(19) => ReadData(19), A(18) => 
                           ReadData(18), A(17) => ReadData(17), A(16) => 
                           ReadData(16), A(15) => ReadData(15), A(14) => 
                           ReadData(14), A(13) => ReadData(13), A(12) => 
                           ReadData(12), A(11) => ReadData(11), A(10) => 
                           ReadData(10), A(9) => ReadData(9), A(8) => 
                           ReadData(8), A(7) => ReadData(7), A(6) => 
                           ReadData(6), A(5) => ReadData(5), A(4) => 
                           ReadData(4), A(3) => ReadData(3), A(2) => 
                           ReadData(2), A(1) => ReadData(1), A(0) => 
                           ReadData(0), B(31) => AluResult(31), B(30) => 
                           AluResult(30), B(29) => AluResult(29), B(28) => 
                           AluResult(28), B(27) => AluResult(27), B(26) => 
                           AluResult(26), B(25) => AluResult(25), B(24) => 
                           AluResult(24), B(23) => AluResult(23), B(22) => 
                           AluResult(22), B(21) => AluResult(21), B(20) => 
                           AluResult(20), B(19) => AluResult(19), B(18) => 
                           AluResult(18), B(17) => AluResult(17), B(16) => 
                           AluResult(16), B(15) => AluResult(15), B(14) => 
                           AluResult(14), B(13) => AluResult(13), B(12) => 
                           AluResult(12), B(11) => AluResult(11), B(10) => 
                           AluResult(10), B(9) => AluResult(9), B(8) => 
                           AluResult(8), B(7) => AluResult(7), B(6) => 
                           AluResult(6), B(5) => AluResult(5), B(4) => 
                           AluResult(4), B(3) => AluResult(3), B(2) => 
                           AluResult(2), B(1) => AluResult(1), B(0) => 
                           AluResult(0), SEL => MemtoReg, Y(31) => 
                           WriteData(31), Y(30) => WriteData(30), Y(29) => 
                           WriteData(29), Y(28) => WriteData(28), Y(27) => 
                           WriteData(27), Y(26) => WriteData(26), Y(25) => 
                           WriteData(25), Y(24) => WriteData(24), Y(23) => 
                           WriteData(23), Y(22) => WriteData(22), Y(21) => 
                           WriteData(21), Y(20) => WriteData(20), Y(19) => 
                           WriteData(19), Y(18) => WriteData(18), Y(17) => 
                           WriteData(17), Y(16) => WriteData(16), Y(15) => 
                           WriteData(15), Y(14) => WriteData(14), Y(13) => 
                           WriteData(13), Y(12) => WriteData(12), Y(11) => 
                           WriteData(11), Y(10) => WriteData(10), Y(9) => 
                           WriteData(9), Y(8) => WriteData(8), Y(7) => 
                           WriteData(7), Y(6) => WriteData(6), Y(5) => 
                           WriteData(5), Y(4) => WriteData(4), Y(3) => 
                           WriteData(3), Y(2) => WriteData(2), Y(1) => 
                           WriteData(1), Y(0) => WriteData(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity memoryUnit_nbit32 is

   port( rst, clk, en_reg, b_op, j_op, jal_op : in std_logic;  alu_out, r2_out,
         PC, lab_b, lab_j, rw_exe, dataout_from_mem : in std_logic_vector (31 
         downto 0);  addr_mem, datain_mem, next_PC, alu_out_mem, rw_mem, 
         data_out : out std_logic_vector (31 downto 0));

end memoryUnit_nbit32;

architecture SYN_struct of memoryUnit_nbit32 is

   component REG_GEN_NBIT32_1
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_2
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_3
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component branch_block_nbit32
      port( branch_op : in std_logic;  cmp_out, PC, label_PC : in 
            std_logic_vector (31 downto 0);  next_PC : out std_logic_vector (31
            downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, branch_pc_31_port, branch_pc_30_port, 
      branch_pc_29_port, branch_pc_28_port, branch_pc_27_port, 
      branch_pc_26_port, branch_pc_25_port, branch_pc_24_port, 
      branch_pc_23_port, branch_pc_22_port, branch_pc_21_port, 
      branch_pc_20_port, branch_pc_19_port, branch_pc_18_port, 
      branch_pc_17_port, branch_pc_16_port, branch_pc_15_port, 
      branch_pc_14_port, branch_pc_13_port, branch_pc_12_port, 
      branch_pc_11_port, branch_pc_10_port, branch_pc_9_port, branch_pc_8_port,
      branch_pc_7_port, branch_pc_6_port, branch_pc_5_port, branch_pc_4_port, 
      branch_pc_3_port, branch_pc_2_port, branch_pc_1_port, branch_pc_0_port, 
      rf_out_31_port, rf_out_30_port, rf_out_29_port, rf_out_28_port, 
      rf_out_27_port, rf_out_26_port, rf_out_25_port, rf_out_24_port, 
      rf_out_23_port, rf_out_22_port, rf_out_21_port, rf_out_20_port, 
      rf_out_19_port, rf_out_18_port, rf_out_17_port, rf_out_16_port, 
      rf_out_15_port, rf_out_14_port, rf_out_13_port, rf_out_12_port, 
      rf_out_11_port, rf_out_10_port, rf_out_9_port, rf_out_8_port, 
      rf_out_7_port, rf_out_6_port, rf_out_5_port, rf_out_4_port, rf_out_3_port
      , rf_out_2_port, rf_out_1_port, rf_out_0_port, rw_out_31_port, 
      rw_out_30_port, rw_out_29_port, rw_out_28_port, rw_out_27_port, 
      rw_out_26_port, rw_out_25_port, rw_out_24_port, rw_out_23_port, 
      rw_out_22_port, rw_out_21_port, rw_out_20_port, rw_out_19_port, 
      rw_out_18_port, rw_out_17_port, rw_out_16_port, rw_out_15_port, 
      rw_out_14_port, rw_out_13_port, rw_out_12_port, rw_out_11_port, 
      rw_out_10_port, rw_out_9_port, rw_out_8_port, rw_out_7_port, 
      rw_out_6_port, rw_out_5_port, rw_out_4_port, rw_out_3_port, rw_out_2_port
      , rw_out_1_port, rw_out_0_port : std_logic;

begin
   addr_mem <= ( alu_out(31), alu_out(30), alu_out(29), alu_out(28), 
      alu_out(27), alu_out(26), alu_out(25), alu_out(24), alu_out(23), 
      alu_out(22), alu_out(21), alu_out(20), alu_out(19), alu_out(18), 
      alu_out(17), alu_out(16), alu_out(15), alu_out(14), alu_out(13), 
      alu_out(12), alu_out(11), alu_out(10), alu_out(9), alu_out(8), alu_out(7)
      , alu_out(6), alu_out(5), alu_out(4), alu_out(3), alu_out(2), alu_out(1),
      alu_out(0) );
   datain_mem <= ( r2_out(31), r2_out(30), r2_out(29), r2_out(28), r2_out(27), 
      r2_out(26), r2_out(25), r2_out(24), r2_out(23), r2_out(22), r2_out(21), 
      r2_out(20), r2_out(19), r2_out(18), r2_out(17), r2_out(16), r2_out(15), 
      r2_out(14), r2_out(13), r2_out(12), r2_out(11), r2_out(10), r2_out(9), 
      r2_out(8), r2_out(7), r2_out(6), r2_out(5), r2_out(4), r2_out(3), 
      r2_out(2), r2_out(1), r2_out(0) );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   br_unit : branch_block_nbit32 port map( branch_op => b_op, cmp_out(31) => 
                           alu_out(31), cmp_out(30) => alu_out(30), cmp_out(29)
                           => alu_out(29), cmp_out(28) => alu_out(28), 
                           cmp_out(27) => alu_out(27), cmp_out(26) => 
                           alu_out(26), cmp_out(25) => alu_out(25), cmp_out(24)
                           => alu_out(24), cmp_out(23) => alu_out(23), 
                           cmp_out(22) => alu_out(22), cmp_out(21) => 
                           alu_out(21), cmp_out(20) => alu_out(20), cmp_out(19)
                           => alu_out(19), cmp_out(18) => alu_out(18), 
                           cmp_out(17) => alu_out(17), cmp_out(16) => 
                           alu_out(16), cmp_out(15) => alu_out(15), cmp_out(14)
                           => alu_out(14), cmp_out(13) => alu_out(13), 
                           cmp_out(12) => alu_out(12), cmp_out(11) => 
                           alu_out(11), cmp_out(10) => alu_out(10), cmp_out(9) 
                           => alu_out(9), cmp_out(8) => alu_out(8), cmp_out(7) 
                           => alu_out(7), cmp_out(6) => alu_out(6), cmp_out(5) 
                           => alu_out(5), cmp_out(4) => alu_out(4), cmp_out(3) 
                           => alu_out(3), cmp_out(2) => alu_out(2), cmp_out(1) 
                           => alu_out(1), cmp_out(0) => alu_out(0), PC(31) => 
                           PC(31), PC(30) => PC(30), PC(29) => PC(29), PC(28) 
                           => PC(28), PC(27) => PC(27), PC(26) => PC(26), 
                           PC(25) => PC(25), PC(24) => PC(24), PC(23) => PC(23)
                           , PC(22) => PC(22), PC(21) => PC(21), PC(20) => 
                           PC(20), PC(19) => PC(19), PC(18) => PC(18), PC(17) 
                           => PC(17), PC(16) => PC(16), PC(15) => PC(15), 
                           PC(14) => PC(14), PC(13) => PC(13), PC(12) => PC(12)
                           , PC(11) => PC(11), PC(10) => PC(10), PC(9) => PC(9)
                           , PC(8) => PC(8), PC(7) => PC(7), PC(6) => PC(6), 
                           PC(5) => PC(5), PC(4) => PC(4), PC(3) => PC(3), 
                           PC(2) => PC(2), PC(1) => PC(1), PC(0) => PC(0), 
                           label_PC(31) => lab_b(31), label_PC(30) => lab_b(30)
                           , label_PC(29) => lab_b(29), label_PC(28) => 
                           lab_b(28), label_PC(27) => lab_b(27), label_PC(26) 
                           => lab_b(26), label_PC(25) => lab_b(25), 
                           label_PC(24) => lab_b(24), label_PC(23) => lab_b(23)
                           , label_PC(22) => lab_b(22), label_PC(21) => 
                           lab_b(21), label_PC(20) => lab_b(20), label_PC(19) 
                           => lab_b(19), label_PC(18) => lab_b(18), 
                           label_PC(17) => lab_b(17), label_PC(16) => lab_b(16)
                           , label_PC(15) => lab_b(15), label_PC(14) => 
                           lab_b(14), label_PC(13) => lab_b(13), label_PC(12) 
                           => lab_b(12), label_PC(11) => lab_b(11), 
                           label_PC(10) => lab_b(10), label_PC(9) => lab_b(9), 
                           label_PC(8) => lab_b(8), label_PC(7) => lab_b(7), 
                           label_PC(6) => lab_b(6), label_PC(5) => lab_b(5), 
                           label_PC(4) => lab_b(4), label_PC(3) => lab_b(3), 
                           label_PC(2) => lab_b(2), label_PC(1) => lab_b(1), 
                           label_PC(0) => lab_b(0), next_PC(31) => 
                           branch_pc_31_port, next_PC(30) => branch_pc_30_port,
                           next_PC(29) => branch_pc_29_port, next_PC(28) => 
                           branch_pc_28_port, next_PC(27) => branch_pc_27_port,
                           next_PC(26) => branch_pc_26_port, next_PC(25) => 
                           branch_pc_25_port, next_PC(24) => branch_pc_24_port,
                           next_PC(23) => branch_pc_23_port, next_PC(22) => 
                           branch_pc_22_port, next_PC(21) => branch_pc_21_port,
                           next_PC(20) => branch_pc_20_port, next_PC(19) => 
                           branch_pc_19_port, next_PC(18) => branch_pc_18_port,
                           next_PC(17) => branch_pc_17_port, next_PC(16) => 
                           branch_pc_16_port, next_PC(15) => branch_pc_15_port,
                           next_PC(14) => branch_pc_14_port, next_PC(13) => 
                           branch_pc_13_port, next_PC(12) => branch_pc_12_port,
                           next_PC(11) => branch_pc_11_port, next_PC(10) => 
                           branch_pc_10_port, next_PC(9) => branch_pc_9_port, 
                           next_PC(8) => branch_pc_8_port, next_PC(7) => 
                           branch_pc_7_port, next_PC(6) => branch_pc_6_port, 
                           next_PC(5) => branch_pc_5_port, next_PC(4) => 
                           branch_pc_4_port, next_PC(3) => branch_pc_3_port, 
                           next_PC(2) => branch_pc_2_port, next_PC(1) => 
                           branch_pc_1_port, next_PC(0) => branch_pc_0_port);
   jmp_unit : MUX21_GENERIC_NBIT32_6 port map( A(31) => branch_pc_31_port, 
                           A(30) => branch_pc_30_port, A(29) => 
                           branch_pc_29_port, A(28) => branch_pc_28_port, A(27)
                           => branch_pc_27_port, A(26) => branch_pc_26_port, 
                           A(25) => branch_pc_25_port, A(24) => 
                           branch_pc_24_port, A(23) => branch_pc_23_port, A(22)
                           => branch_pc_22_port, A(21) => branch_pc_21_port, 
                           A(20) => branch_pc_20_port, A(19) => 
                           branch_pc_19_port, A(18) => branch_pc_18_port, A(17)
                           => branch_pc_17_port, A(16) => branch_pc_16_port, 
                           A(15) => branch_pc_15_port, A(14) => 
                           branch_pc_14_port, A(13) => branch_pc_13_port, A(12)
                           => branch_pc_12_port, A(11) => branch_pc_11_port, 
                           A(10) => branch_pc_10_port, A(9) => branch_pc_9_port
                           , A(8) => branch_pc_8_port, A(7) => branch_pc_7_port
                           , A(6) => branch_pc_6_port, A(5) => branch_pc_5_port
                           , A(4) => branch_pc_4_port, A(3) => branch_pc_3_port
                           , A(2) => branch_pc_2_port, A(1) => branch_pc_1_port
                           , A(0) => branch_pc_0_port, B(31) => lab_j(31), 
                           B(30) => lab_j(30), B(29) => lab_j(29), B(28) => 
                           lab_j(28), B(27) => lab_j(27), B(26) => lab_j(26), 
                           B(25) => lab_j(25), B(24) => lab_j(24), B(23) => 
                           lab_j(23), B(22) => lab_j(22), B(21) => lab_j(21), 
                           B(20) => lab_j(20), B(19) => lab_j(19), B(18) => 
                           lab_j(18), B(17) => lab_j(17), B(16) => lab_j(16), 
                           B(15) => lab_j(15), B(14) => lab_j(14), B(13) => 
                           lab_j(13), B(12) => lab_j(12), B(11) => lab_j(11), 
                           B(10) => lab_j(10), B(9) => lab_j(9), B(8) => 
                           lab_j(8), B(7) => lab_j(7), B(6) => lab_j(6), B(5) 
                           => lab_j(5), B(4) => lab_j(4), B(3) => lab_j(3), 
                           B(2) => lab_j(2), B(1) => lab_j(1), B(0) => lab_j(0)
                           , SEL => j_op, Y(31) => next_PC(31), Y(30) => 
                           next_PC(30), Y(29) => next_PC(29), Y(28) => 
                           next_PC(28), Y(27) => next_PC(27), Y(26) => 
                           next_PC(26), Y(25) => next_PC(25), Y(24) => 
                           next_PC(24), Y(23) => next_PC(23), Y(22) => 
                           next_PC(22), Y(21) => next_PC(21), Y(20) => 
                           next_PC(20), Y(19) => next_PC(19), Y(18) => 
                           next_PC(18), Y(17) => next_PC(17), Y(16) => 
                           next_PC(16), Y(15) => next_PC(15), Y(14) => 
                           next_PC(14), Y(13) => next_PC(13), Y(12) => 
                           next_PC(12), Y(11) => next_PC(11), Y(10) => 
                           next_PC(10), Y(9) => next_PC(9), Y(8) => next_PC(8),
                           Y(7) => next_PC(7), Y(6) => next_PC(6), Y(5) => 
                           next_PC(5), Y(4) => next_PC(4), Y(3) => next_PC(3), 
                           Y(2) => next_PC(2), Y(1) => next_PC(1), Y(0) => 
                           next_PC(0));
   mux_jal_pc : MUX21_GENERIC_NBIT32_5 port map( A(31) => dataout_from_mem(31),
                           A(30) => dataout_from_mem(30), A(29) => 
                           dataout_from_mem(29), A(28) => dataout_from_mem(28),
                           A(27) => dataout_from_mem(27), A(26) => 
                           dataout_from_mem(26), A(25) => dataout_from_mem(25),
                           A(24) => dataout_from_mem(24), A(23) => 
                           dataout_from_mem(23), A(22) => dataout_from_mem(22),
                           A(21) => dataout_from_mem(21), A(20) => 
                           dataout_from_mem(20), A(19) => dataout_from_mem(19),
                           A(18) => dataout_from_mem(18), A(17) => 
                           dataout_from_mem(17), A(16) => dataout_from_mem(16),
                           A(15) => dataout_from_mem(15), A(14) => 
                           dataout_from_mem(14), A(13) => dataout_from_mem(13),
                           A(12) => dataout_from_mem(12), A(11) => 
                           dataout_from_mem(11), A(10) => dataout_from_mem(10),
                           A(9) => dataout_from_mem(9), A(8) => 
                           dataout_from_mem(8), A(7) => dataout_from_mem(7), 
                           A(6) => dataout_from_mem(6), A(5) => 
                           dataout_from_mem(5), A(4) => dataout_from_mem(4), 
                           A(3) => dataout_from_mem(3), A(2) => 
                           dataout_from_mem(2), A(1) => dataout_from_mem(1), 
                           A(0) => dataout_from_mem(0), B(31) => PC(31), B(30) 
                           => PC(30), B(29) => PC(29), B(28) => PC(28), B(27) 
                           => PC(27), B(26) => PC(26), B(25) => PC(25), B(24) 
                           => PC(24), B(23) => PC(23), B(22) => PC(22), B(21) 
                           => PC(21), B(20) => PC(20), B(19) => PC(19), B(18) 
                           => PC(18), B(17) => PC(17), B(16) => PC(16), B(15) 
                           => PC(15), B(14) => PC(14), B(13) => PC(13), B(12) 
                           => PC(12), B(11) => PC(11), B(10) => PC(10), B(9) =>
                           PC(9), B(8) => PC(8), B(7) => PC(7), B(6) => PC(6), 
                           B(5) => PC(5), B(4) => PC(4), B(3) => PC(3), B(2) =>
                           PC(2), B(1) => PC(1), B(0) => PC(0), SEL => jal_op, 
                           Y(31) => rf_out_31_port, Y(30) => rf_out_30_port, 
                           Y(29) => rf_out_29_port, Y(28) => rf_out_28_port, 
                           Y(27) => rf_out_27_port, Y(26) => rf_out_26_port, 
                           Y(25) => rf_out_25_port, Y(24) => rf_out_24_port, 
                           Y(23) => rf_out_23_port, Y(22) => rf_out_22_port, 
                           Y(21) => rf_out_21_port, Y(20) => rf_out_20_port, 
                           Y(19) => rf_out_19_port, Y(18) => rf_out_18_port, 
                           Y(17) => rf_out_17_port, Y(16) => rf_out_16_port, 
                           Y(15) => rf_out_15_port, Y(14) => rf_out_14_port, 
                           Y(13) => rf_out_13_port, Y(12) => rf_out_12_port, 
                           Y(11) => rf_out_11_port, Y(10) => rf_out_10_port, 
                           Y(9) => rf_out_9_port, Y(8) => rf_out_8_port, Y(7) 
                           => rf_out_7_port, Y(6) => rf_out_6_port, Y(5) => 
                           rf_out_5_port, Y(4) => rf_out_4_port, Y(3) => 
                           rf_out_3_port, Y(2) => rf_out_2_port, Y(1) => 
                           rf_out_1_port, Y(0) => rf_out_0_port);
   mux_jal_r31 : MUX21_GENERIC_NBIT32_4 port map( A(31) => rw_exe(31), A(30) =>
                           rw_exe(30), A(29) => rw_exe(29), A(28) => rw_exe(28)
                           , A(27) => rw_exe(27), A(26) => rw_exe(26), A(25) =>
                           rw_exe(25), A(24) => rw_exe(24), A(23) => rw_exe(23)
                           , A(22) => rw_exe(22), A(21) => rw_exe(21), A(20) =>
                           rw_exe(20), A(19) => rw_exe(19), A(18) => rw_exe(18)
                           , A(17) => rw_exe(17), A(16) => rw_exe(16), A(15) =>
                           rw_exe(15), A(14) => rw_exe(14), A(13) => rw_exe(13)
                           , A(12) => rw_exe(12), A(11) => rw_exe(11), A(10) =>
                           rw_exe(10), A(9) => rw_exe(9), A(8) => rw_exe(8), 
                           A(7) => rw_exe(7), A(6) => rw_exe(6), A(5) => 
                           rw_exe(5), A(4) => rw_exe(4), A(3) => rw_exe(3), 
                           A(2) => rw_exe(2), A(1) => rw_exe(1), A(0) => 
                           rw_exe(0), B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic1_port, B(3) => X_Logic1_port, B(2) => 
                           X_Logic1_port, B(1) => X_Logic1_port, B(0) => 
                           X_Logic1_port, SEL => jal_op, Y(31) => 
                           rw_out_31_port, Y(30) => rw_out_30_port, Y(29) => 
                           rw_out_29_port, Y(28) => rw_out_28_port, Y(27) => 
                           rw_out_27_port, Y(26) => rw_out_26_port, Y(25) => 
                           rw_out_25_port, Y(24) => rw_out_24_port, Y(23) => 
                           rw_out_23_port, Y(22) => rw_out_22_port, Y(21) => 
                           rw_out_21_port, Y(20) => rw_out_20_port, Y(19) => 
                           rw_out_19_port, Y(18) => rw_out_18_port, Y(17) => 
                           rw_out_17_port, Y(16) => rw_out_16_port, Y(15) => 
                           rw_out_15_port, Y(14) => rw_out_14_port, Y(13) => 
                           rw_out_13_port, Y(12) => rw_out_12_port, Y(11) => 
                           rw_out_11_port, Y(10) => rw_out_10_port, Y(9) => 
                           rw_out_9_port, Y(8) => rw_out_8_port, Y(7) => 
                           rw_out_7_port, Y(6) => rw_out_6_port, Y(5) => 
                           rw_out_5_port, Y(4) => rw_out_4_port, Y(3) => 
                           rw_out_3_port, Y(2) => rw_out_2_port, Y(1) => 
                           rw_out_1_port, Y(0) => rw_out_0_port);
   mem_reg : REG_GEN_NBIT32_3 port map( D(31) => rf_out_31_port, D(30) => 
                           rf_out_30_port, D(29) => rf_out_29_port, D(28) => 
                           rf_out_28_port, D(27) => rf_out_27_port, D(26) => 
                           rf_out_26_port, D(25) => rf_out_25_port, D(24) => 
                           rf_out_24_port, D(23) => rf_out_23_port, D(22) => 
                           rf_out_22_port, D(21) => rf_out_21_port, D(20) => 
                           rf_out_20_port, D(19) => rf_out_19_port, D(18) => 
                           rf_out_18_port, D(17) => rf_out_17_port, D(16) => 
                           rf_out_16_port, D(15) => rf_out_15_port, D(14) => 
                           rf_out_14_port, D(13) => rf_out_13_port, D(12) => 
                           rf_out_12_port, D(11) => rf_out_11_port, D(10) => 
                           rf_out_10_port, D(9) => rf_out_9_port, D(8) => 
                           rf_out_8_port, D(7) => rf_out_7_port, D(6) => 
                           rf_out_6_port, D(5) => rf_out_5_port, D(4) => 
                           rf_out_4_port, D(3) => rf_out_3_port, D(2) => 
                           rf_out_2_port, D(1) => rf_out_1_port, D(0) => 
                           rf_out_0_port, CK => clk, Enable_n => en_reg, 
                           RESET_n => rst, Q(31) => data_out(31), Q(30) => 
                           data_out(30), Q(29) => data_out(29), Q(28) => 
                           data_out(28), Q(27) => data_out(27), Q(26) => 
                           data_out(26), Q(25) => data_out(25), Q(24) => 
                           data_out(24), Q(23) => data_out(23), Q(22) => 
                           data_out(22), Q(21) => data_out(21), Q(20) => 
                           data_out(20), Q(19) => data_out(19), Q(18) => 
                           data_out(18), Q(17) => data_out(17), Q(16) => 
                           data_out(16), Q(15) => data_out(15), Q(14) => 
                           data_out(14), Q(13) => data_out(13), Q(12) => 
                           data_out(12), Q(11) => data_out(11), Q(10) => 
                           data_out(10), Q(9) => data_out(9), Q(8) => 
                           data_out(8), Q(7) => data_out(7), Q(6) => 
                           data_out(6), Q(5) => data_out(5), Q(4) => 
                           data_out(4), Q(3) => data_out(3), Q(2) => 
                           data_out(2), Q(1) => data_out(1), Q(0) => 
                           data_out(0));
   rw_reg : REG_GEN_NBIT32_2 port map( D(31) => rw_out_31_port, D(30) => 
                           rw_out_30_port, D(29) => rw_out_29_port, D(28) => 
                           rw_out_28_port, D(27) => rw_out_27_port, D(26) => 
                           rw_out_26_port, D(25) => rw_out_25_port, D(24) => 
                           rw_out_24_port, D(23) => rw_out_23_port, D(22) => 
                           rw_out_22_port, D(21) => rw_out_21_port, D(20) => 
                           rw_out_20_port, D(19) => rw_out_19_port, D(18) => 
                           rw_out_18_port, D(17) => rw_out_17_port, D(16) => 
                           rw_out_16_port, D(15) => rw_out_15_port, D(14) => 
                           rw_out_14_port, D(13) => rw_out_13_port, D(12) => 
                           rw_out_12_port, D(11) => rw_out_11_port, D(10) => 
                           rw_out_10_port, D(9) => rw_out_9_port, D(8) => 
                           rw_out_8_port, D(7) => rw_out_7_port, D(6) => 
                           rw_out_6_port, D(5) => rw_out_5_port, D(4) => 
                           rw_out_4_port, D(3) => rw_out_3_port, D(2) => 
                           rw_out_2_port, D(1) => rw_out_1_port, D(0) => 
                           rw_out_0_port, CK => clk, Enable_n => en_reg, 
                           RESET_n => rst, Q(31) => rw_mem(31), Q(30) => 
                           rw_mem(30), Q(29) => rw_mem(29), Q(28) => rw_mem(28)
                           , Q(27) => rw_mem(27), Q(26) => rw_mem(26), Q(25) =>
                           rw_mem(25), Q(24) => rw_mem(24), Q(23) => rw_mem(23)
                           , Q(22) => rw_mem(22), Q(21) => rw_mem(21), Q(20) =>
                           rw_mem(20), Q(19) => rw_mem(19), Q(18) => rw_mem(18)
                           , Q(17) => rw_mem(17), Q(16) => rw_mem(16), Q(15) =>
                           rw_mem(15), Q(14) => rw_mem(14), Q(13) => rw_mem(13)
                           , Q(12) => rw_mem(12), Q(11) => rw_mem(11), Q(10) =>
                           rw_mem(10), Q(9) => rw_mem(9), Q(8) => rw_mem(8), 
                           Q(7) => rw_mem(7), Q(6) => rw_mem(6), Q(5) => 
                           rw_mem(5), Q(4) => rw_mem(4), Q(3) => rw_mem(3), 
                           Q(2) => rw_mem(2), Q(1) => rw_mem(1), Q(0) => 
                           rw_mem(0));
   alu_reg : REG_GEN_NBIT32_1 port map( D(31) => alu_out(31), D(30) => 
                           alu_out(30), D(29) => alu_out(29), D(28) => 
                           alu_out(28), D(27) => alu_out(27), D(26) => 
                           alu_out(26), D(25) => alu_out(25), D(24) => 
                           alu_out(24), D(23) => alu_out(23), D(22) => 
                           alu_out(22), D(21) => alu_out(21), D(20) => 
                           alu_out(20), D(19) => alu_out(19), D(18) => 
                           alu_out(18), D(17) => alu_out(17), D(16) => 
                           alu_out(16), D(15) => alu_out(15), D(14) => 
                           alu_out(14), D(13) => alu_out(13), D(12) => 
                           alu_out(12), D(11) => alu_out(11), D(10) => 
                           alu_out(10), D(9) => alu_out(9), D(8) => alu_out(8),
                           D(7) => alu_out(7), D(6) => alu_out(6), D(5) => 
                           alu_out(5), D(4) => alu_out(4), D(3) => alu_out(3), 
                           D(2) => alu_out(2), D(1) => alu_out(1), D(0) => 
                           alu_out(0), CK => clk, Enable_n => en_reg, RESET_n 
                           => rst, Q(31) => alu_out_mem(31), Q(30) => 
                           alu_out_mem(30), Q(29) => alu_out_mem(29), Q(28) => 
                           alu_out_mem(28), Q(27) => alu_out_mem(27), Q(26) => 
                           alu_out_mem(26), Q(25) => alu_out_mem(25), Q(24) => 
                           alu_out_mem(24), Q(23) => alu_out_mem(23), Q(22) => 
                           alu_out_mem(22), Q(21) => alu_out_mem(21), Q(20) => 
                           alu_out_mem(20), Q(19) => alu_out_mem(19), Q(18) => 
                           alu_out_mem(18), Q(17) => alu_out_mem(17), Q(16) => 
                           alu_out_mem(16), Q(15) => alu_out_mem(15), Q(14) => 
                           alu_out_mem(14), Q(13) => alu_out_mem(13), Q(12) => 
                           alu_out_mem(12), Q(11) => alu_out_mem(11), Q(10) => 
                           alu_out_mem(10), Q(9) => alu_out_mem(9), Q(8) => 
                           alu_out_mem(8), Q(7) => alu_out_mem(7), Q(6) => 
                           alu_out_mem(6), Q(5) => alu_out_mem(5), Q(4) => 
                           alu_out_mem(4), Q(3) => alu_out_mem(3), Q(2) => 
                           alu_out_mem(2), Q(1) => alu_out_mem(1), Q(0) => 
                           alu_out_mem(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity executionUnit_nbit32 is

   port( r1, r2, imm, j_lab, pc, RW_R, RW_I : in std_logic_vector (31 downto 0)
         ;  s2, s3, rst, clk, en_reg : in std_logic;  alu_sel : in 
         std_logic_vector (3 downto 0);  alu_out, alu_fw_out, r2_out, b_lab_out
         , pc_exe_out, rw_exe, j_lab_out : out std_logic_vector (31 downto 0));

end executionUnit_nbit32;

architecture SYN_struct of executionUnit_nbit32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component REG_GEN_NBIT32_4
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_5
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_6
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_7
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component P4_ADDER_NBIT32_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component P4_ADDER_NBIT32_NBIT_PER_BLOCK4_3
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_8
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_9
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component alu
      port( data_in1, data_in2 : in std_logic_vector (31 downto 0);  op_sel : 
            in std_logic_vector (3 downto 0);  data_out : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_7
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_8
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, alu_fw_out_31_port, alu_fw_out_30_port, 
      alu_fw_out_29_port, alu_fw_out_28_port, alu_fw_out_27_port, 
      alu_fw_out_26_port, alu_fw_out_25_port, alu_fw_out_24_port, 
      alu_fw_out_23_port, alu_fw_out_22_port, alu_fw_out_21_port, 
      alu_fw_out_20_port, alu_fw_out_19_port, alu_fw_out_18_port, 
      alu_fw_out_17_port, alu_fw_out_16_port, alu_fw_out_15_port, 
      alu_fw_out_14_port, alu_fw_out_13_port, alu_fw_out_12_port, 
      alu_fw_out_11_port, alu_fw_out_10_port, alu_fw_out_9_port, 
      alu_fw_out_8_port, alu_fw_out_7_port, alu_fw_out_6_port, 
      alu_fw_out_5_port, alu_fw_out_4_port, alu_fw_out_3_port, 
      alu_fw_out_2_port, alu_fw_out_1_port, alu_fw_out_0_port, mux_out_31_port,
      mux_out_30_port, mux_out_29_port, mux_out_28_port, mux_out_27_port, 
      mux_out_26_port, mux_out_25_port, mux_out_24_port, mux_out_23_port, 
      mux_out_22_port, mux_out_21_port, mux_out_20_port, mux_out_19_port, 
      mux_out_18_port, mux_out_17_port, mux_out_16_port, mux_out_15_port, 
      mux_out_14_port, mux_out_13_port, mux_out_12_port, mux_out_11_port, 
      mux_out_10_port, mux_out_9_port, mux_out_8_port, mux_out_7_port, 
      mux_out_6_port, mux_out_5_port, mux_out_4_port, mux_out_3_port, 
      mux_out_2_port, mux_out_1_port, mux_out_0_port, rw_s_31_port, 
      rw_s_30_port, rw_s_29_port, rw_s_28_port, rw_s_27_port, rw_s_26_port, 
      rw_s_25_port, rw_s_24_port, rw_s_23_port, rw_s_22_port, rw_s_21_port, 
      rw_s_20_port, rw_s_19_port, rw_s_18_port, rw_s_17_port, rw_s_16_port, 
      rw_s_15_port, rw_s_14_port, rw_s_13_port, rw_s_12_port, rw_s_11_port, 
      rw_s_10_port, rw_s_9_port, rw_s_8_port, rw_s_7_port, rw_s_6_port, 
      rw_s_5_port, rw_s_4_port, rw_s_3_port, rw_s_2_port, rw_s_1_port, 
      rw_s_0_port, pc_b_31_port, pc_b_30_port, pc_b_29_port, pc_b_28_port, 
      pc_b_27_port, pc_b_26_port, pc_b_25_port, pc_b_24_port, pc_b_23_port, 
      pc_b_22_port, pc_b_21_port, pc_b_20_port, pc_b_19_port, pc_b_18_port, 
      pc_b_17_port, pc_b_16_port, pc_b_15_port, pc_b_14_port, pc_b_13_port, 
      pc_b_12_port, pc_b_11_port, pc_b_10_port, pc_b_9_port, pc_b_8_port, 
      pc_b_7_port, pc_b_6_port, pc_b_5_port, pc_b_4_port, pc_b_3_port, 
      pc_b_2_port, pc_b_1_port, pc_b_0_port, pc_j_31_port, pc_j_30_port, 
      pc_j_29_port, pc_j_28_port, pc_j_27_port, pc_j_26_port, pc_j_25_port, 
      pc_j_24_port, pc_j_23_port, pc_j_22_port, pc_j_21_port, pc_j_20_port, 
      pc_j_19_port, pc_j_18_port, pc_j_17_port, pc_j_16_port, pc_j_15_port, 
      pc_j_14_port, pc_j_13_port, pc_j_12_port, pc_j_11_port, pc_j_10_port, 
      pc_j_9_port, pc_j_8_port, pc_j_7_port, pc_j_6_port, pc_j_5_port, 
      pc_j_4_port, pc_j_3_port, pc_j_2_port, pc_j_1_port, pc_j_0_port, n1, n2, 
      n_1200, n_1201 : std_logic;

begin
   alu_fw_out <= ( alu_fw_out_31_port, alu_fw_out_30_port, alu_fw_out_29_port, 
      alu_fw_out_28_port, alu_fw_out_27_port, alu_fw_out_26_port, 
      alu_fw_out_25_port, alu_fw_out_24_port, alu_fw_out_23_port, 
      alu_fw_out_22_port, alu_fw_out_21_port, alu_fw_out_20_port, 
      alu_fw_out_19_port, alu_fw_out_18_port, alu_fw_out_17_port, 
      alu_fw_out_16_port, alu_fw_out_15_port, alu_fw_out_14_port, 
      alu_fw_out_13_port, alu_fw_out_12_port, alu_fw_out_11_port, 
      alu_fw_out_10_port, alu_fw_out_9_port, alu_fw_out_8_port, 
      alu_fw_out_7_port, alu_fw_out_6_port, alu_fw_out_5_port, 
      alu_fw_out_4_port, alu_fw_out_3_port, alu_fw_out_2_port, 
      alu_fw_out_1_port, alu_fw_out_0_port );
   
   X_Logic0_port <= '0';
   lo_mux : MUX21_GENERIC_NBIT32_8 port map( A(31) => r2(31), A(30) => r2(30), 
                           A(29) => r2(29), A(28) => r2(28), A(27) => r2(27), 
                           A(26) => r2(26), A(25) => r2(25), A(24) => r2(24), 
                           A(23) => r2(23), A(22) => r2(22), A(21) => r2(21), 
                           A(20) => r2(20), A(19) => r2(19), A(18) => r2(18), 
                           A(17) => r2(17), A(16) => r2(16), A(15) => r2(15), 
                           A(14) => r2(14), A(13) => r2(13), A(12) => r2(12), 
                           A(11) => r2(11), A(10) => r2(10), A(9) => r2(9), 
                           A(8) => r2(8), A(7) => r2(7), A(6) => r2(6), A(5) =>
                           r2(5), A(4) => r2(4), A(3) => r2(3), A(2) => r2(2), 
                           A(1) => r2(1), A(0) => r2(0), B(31) => imm(31), 
                           B(30) => imm(30), B(29) => imm(29), B(28) => imm(28)
                           , B(27) => imm(27), B(26) => imm(26), B(25) => 
                           imm(25), B(24) => imm(24), B(23) => imm(23), B(22) 
                           => imm(22), B(21) => imm(21), B(20) => imm(20), 
                           B(19) => imm(19), B(18) => imm(18), B(17) => imm(17)
                           , B(16) => imm(16), B(15) => imm(15), B(14) => 
                           imm(14), B(13) => imm(13), B(12) => imm(12), B(11) 
                           => imm(11), B(10) => imm(10), B(9) => imm(9), B(8) 
                           => imm(8), B(7) => imm(7), B(6) => imm(6), B(5) => 
                           imm(5), B(4) => imm(4), B(3) => imm(3), B(2) => 
                           imm(2), B(1) => imm(1), B(0) => imm(0), SEL => s2, 
                           Y(31) => mux_out_31_port, Y(30) => mux_out_30_port, 
                           Y(29) => mux_out_29_port, Y(28) => mux_out_28_port, 
                           Y(27) => mux_out_27_port, Y(26) => mux_out_26_port, 
                           Y(25) => mux_out_25_port, Y(24) => mux_out_24_port, 
                           Y(23) => mux_out_23_port, Y(22) => mux_out_22_port, 
                           Y(21) => mux_out_21_port, Y(20) => mux_out_20_port, 
                           Y(19) => mux_out_19_port, Y(18) => mux_out_18_port, 
                           Y(17) => mux_out_17_port, Y(16) => mux_out_16_port, 
                           Y(15) => mux_out_15_port, Y(14) => mux_out_14_port, 
                           Y(13) => mux_out_13_port, Y(12) => mux_out_12_port, 
                           Y(11) => mux_out_11_port, Y(10) => mux_out_10_port, 
                           Y(9) => mux_out_9_port, Y(8) => mux_out_8_port, Y(7)
                           => mux_out_7_port, Y(6) => mux_out_6_port, Y(5) => 
                           mux_out_5_port, Y(4) => mux_out_4_port, Y(3) => 
                           mux_out_3_port, Y(2) => mux_out_2_port, Y(1) => 
                           mux_out_1_port, Y(0) => mux_out_0_port);
   RW_mux : MUX21_GENERIC_NBIT32_7 port map( A(31) => RW_R(31), A(30) => 
                           RW_R(30), A(29) => RW_R(29), A(28) => RW_R(28), 
                           A(27) => RW_R(27), A(26) => RW_R(26), A(25) => 
                           RW_R(25), A(24) => RW_R(24), A(23) => RW_R(23), 
                           A(22) => RW_R(22), A(21) => RW_R(21), A(20) => 
                           RW_R(20), A(19) => RW_R(19), A(18) => RW_R(18), 
                           A(17) => RW_R(17), A(16) => RW_R(16), A(15) => 
                           RW_R(15), A(14) => RW_R(14), A(13) => RW_R(13), 
                           A(12) => RW_R(12), A(11) => RW_R(11), A(10) => 
                           RW_R(10), A(9) => RW_R(9), A(8) => RW_R(8), A(7) => 
                           RW_R(7), A(6) => RW_R(6), A(5) => RW_R(5), A(4) => 
                           RW_R(4), A(3) => RW_R(3), A(2) => RW_R(2), A(1) => 
                           RW_R(1), A(0) => RW_R(0), B(31) => RW_I(31), B(30) 
                           => RW_I(30), B(29) => RW_I(29), B(28) => RW_I(28), 
                           B(27) => RW_I(27), B(26) => RW_I(26), B(25) => 
                           RW_I(25), B(24) => RW_I(24), B(23) => RW_I(23), 
                           B(22) => RW_I(22), B(21) => RW_I(21), B(20) => 
                           RW_I(20), B(19) => RW_I(19), B(18) => RW_I(18), 
                           B(17) => RW_I(17), B(16) => RW_I(16), B(15) => 
                           RW_I(15), B(14) => RW_I(14), B(13) => RW_I(13), 
                           B(12) => RW_I(12), B(11) => RW_I(11), B(10) => 
                           RW_I(10), B(9) => RW_I(9), B(8) => RW_I(8), B(7) => 
                           RW_I(7), B(6) => RW_I(6), B(5) => RW_I(5), B(4) => 
                           RW_I(4), B(3) => RW_I(3), B(2) => RW_I(2), B(1) => 
                           RW_I(1), B(0) => RW_I(0), SEL => s3, Y(31) => 
                           rw_s_31_port, Y(30) => rw_s_30_port, Y(29) => 
                           rw_s_29_port, Y(28) => rw_s_28_port, Y(27) => 
                           rw_s_27_port, Y(26) => rw_s_26_port, Y(25) => 
                           rw_s_25_port, Y(24) => rw_s_24_port, Y(23) => 
                           rw_s_23_port, Y(22) => rw_s_22_port, Y(21) => 
                           rw_s_21_port, Y(20) => rw_s_20_port, Y(19) => 
                           rw_s_19_port, Y(18) => rw_s_18_port, Y(17) => 
                           rw_s_17_port, Y(16) => rw_s_16_port, Y(15) => 
                           rw_s_15_port, Y(14) => rw_s_14_port, Y(13) => 
                           rw_s_13_port, Y(12) => rw_s_12_port, Y(11) => 
                           rw_s_11_port, Y(10) => rw_s_10_port, Y(9) => 
                           rw_s_9_port, Y(8) => rw_s_8_port, Y(7) => 
                           rw_s_7_port, Y(6) => rw_s_6_port, Y(5) => 
                           rw_s_5_port, Y(4) => rw_s_4_port, Y(3) => 
                           rw_s_3_port, Y(2) => rw_s_2_port, Y(1) => 
                           rw_s_1_port, Y(0) => rw_s_0_port);
   alu_dut : alu port map( data_in1(31) => r1(31), data_in1(30) => r1(30), 
                           data_in1(29) => r1(29), data_in1(28) => r1(28), 
                           data_in1(27) => r1(27), data_in1(26) => r1(26), 
                           data_in1(25) => n1, data_in1(24) => r1(24), 
                           data_in1(23) => r1(23), data_in1(22) => r1(22), 
                           data_in1(21) => r1(21), data_in1(20) => r1(20), 
                           data_in1(19) => r1(19), data_in1(18) => r1(18), 
                           data_in1(17) => r1(17), data_in1(16) => r1(16), 
                           data_in1(15) => r1(15), data_in1(14) => r1(14), 
                           data_in1(13) => r1(13), data_in1(12) => r1(12), 
                           data_in1(11) => r1(11), data_in1(10) => r1(10), 
                           data_in1(9) => r1(9), data_in1(8) => r1(8), 
                           data_in1(7) => r1(7), data_in1(6) => r1(6), 
                           data_in1(5) => r1(5), data_in1(4) => r1(4), 
                           data_in1(3) => r1(3), data_in1(2) => r1(2), 
                           data_in1(1) => r1(1), data_in1(0) => r1(0), 
                           data_in2(31) => mux_out_31_port, data_in2(30) => 
                           mux_out_30_port, data_in2(29) => mux_out_29_port, 
                           data_in2(28) => mux_out_28_port, data_in2(27) => 
                           mux_out_27_port, data_in2(26) => mux_out_26_port, 
                           data_in2(25) => mux_out_25_port, data_in2(24) => 
                           mux_out_24_port, data_in2(23) => mux_out_23_port, 
                           data_in2(22) => mux_out_22_port, data_in2(21) => 
                           mux_out_21_port, data_in2(20) => mux_out_20_port, 
                           data_in2(19) => mux_out_19_port, data_in2(18) => 
                           mux_out_18_port, data_in2(17) => mux_out_17_port, 
                           data_in2(16) => mux_out_16_port, data_in2(15) => 
                           mux_out_15_port, data_in2(14) => mux_out_14_port, 
                           data_in2(13) => mux_out_13_port, data_in2(12) => 
                           mux_out_12_port, data_in2(11) => mux_out_11_port, 
                           data_in2(10) => mux_out_10_port, data_in2(9) => 
                           mux_out_9_port, data_in2(8) => mux_out_8_port, 
                           data_in2(7) => mux_out_7_port, data_in2(6) => 
                           mux_out_6_port, data_in2(5) => mux_out_5_port, 
                           data_in2(4) => mux_out_4_port, data_in2(3) => 
                           mux_out_3_port, data_in2(2) => mux_out_2_port, 
                           data_in2(1) => mux_out_1_port, data_in2(0) => 
                           mux_out_0_port, op_sel(3) => alu_sel(3), op_sel(2) 
                           => alu_sel(2), op_sel(1) => alu_sel(1), op_sel(0) =>
                           alu_sel(0), data_out(31) => alu_fw_out_31_port, 
                           data_out(30) => alu_fw_out_30_port, data_out(29) => 
                           alu_fw_out_29_port, data_out(28) => 
                           alu_fw_out_28_port, data_out(27) => 
                           alu_fw_out_27_port, data_out(26) => 
                           alu_fw_out_26_port, data_out(25) => 
                           alu_fw_out_25_port, data_out(24) => 
                           alu_fw_out_24_port, data_out(23) => 
                           alu_fw_out_23_port, data_out(22) => 
                           alu_fw_out_22_port, data_out(21) => 
                           alu_fw_out_21_port, data_out(20) => 
                           alu_fw_out_20_port, data_out(19) => 
                           alu_fw_out_19_port, data_out(18) => 
                           alu_fw_out_18_port, data_out(17) => 
                           alu_fw_out_17_port, data_out(16) => 
                           alu_fw_out_16_port, data_out(15) => 
                           alu_fw_out_15_port, data_out(14) => 
                           alu_fw_out_14_port, data_out(13) => 
                           alu_fw_out_13_port, data_out(12) => 
                           alu_fw_out_12_port, data_out(11) => 
                           alu_fw_out_11_port, data_out(10) => 
                           alu_fw_out_10_port, data_out(9) => alu_fw_out_9_port
                           , data_out(8) => alu_fw_out_8_port, data_out(7) => 
                           alu_fw_out_7_port, data_out(6) => alu_fw_out_6_port,
                           data_out(5) => alu_fw_out_5_port, data_out(4) => 
                           alu_fw_out_4_port, data_out(3) => alu_fw_out_3_port,
                           data_out(2) => alu_fw_out_2_port, data_out(1) => 
                           alu_fw_out_1_port, data_out(0) => alu_fw_out_0_port)
                           ;
   reg_alu : REG_GEN_NBIT32_9 port map( D(31) => alu_fw_out_31_port, D(30) => 
                           alu_fw_out_30_port, D(29) => alu_fw_out_29_port, 
                           D(28) => alu_fw_out_28_port, D(27) => 
                           alu_fw_out_27_port, D(26) => alu_fw_out_26_port, 
                           D(25) => alu_fw_out_25_port, D(24) => 
                           alu_fw_out_24_port, D(23) => alu_fw_out_23_port, 
                           D(22) => alu_fw_out_22_port, D(21) => 
                           alu_fw_out_21_port, D(20) => alu_fw_out_20_port, 
                           D(19) => alu_fw_out_19_port, D(18) => 
                           alu_fw_out_18_port, D(17) => alu_fw_out_17_port, 
                           D(16) => alu_fw_out_16_port, D(15) => 
                           alu_fw_out_15_port, D(14) => alu_fw_out_14_port, 
                           D(13) => alu_fw_out_13_port, D(12) => 
                           alu_fw_out_12_port, D(11) => alu_fw_out_11_port, 
                           D(10) => alu_fw_out_10_port, D(9) => 
                           alu_fw_out_9_port, D(8) => alu_fw_out_8_port, D(7) 
                           => alu_fw_out_7_port, D(6) => alu_fw_out_6_port, 
                           D(5) => alu_fw_out_5_port, D(4) => alu_fw_out_4_port
                           , D(3) => alu_fw_out_3_port, D(2) => 
                           alu_fw_out_2_port, D(1) => alu_fw_out_1_port, D(0) 
                           => alu_fw_out_0_port, CK => clk, Enable_n => n2, 
                           RESET_n => rst, Q(31) => alu_out(31), Q(30) => 
                           alu_out(30), Q(29) => alu_out(29), Q(28) => 
                           alu_out(28), Q(27) => alu_out(27), Q(26) => 
                           alu_out(26), Q(25) => alu_out(25), Q(24) => 
                           alu_out(24), Q(23) => alu_out(23), Q(22) => 
                           alu_out(22), Q(21) => alu_out(21), Q(20) => 
                           alu_out(20), Q(19) => alu_out(19), Q(18) => 
                           alu_out(18), Q(17) => alu_out(17), Q(16) => 
                           alu_out(16), Q(15) => alu_out(15), Q(14) => 
                           alu_out(14), Q(13) => alu_out(13), Q(12) => 
                           alu_out(12), Q(11) => alu_out(11), Q(10) => 
                           alu_out(10), Q(9) => alu_out(9), Q(8) => alu_out(8),
                           Q(7) => alu_out(7), Q(6) => alu_out(6), Q(5) => 
                           alu_out(5), Q(4) => alu_out(4), Q(3) => alu_out(3), 
                           Q(2) => alu_out(2), Q(1) => alu_out(1), Q(0) => 
                           alu_out(0));
   ls_reg : REG_GEN_NBIT32_8 port map( D(31) => r2(31), D(30) => r2(30), D(29) 
                           => r2(29), D(28) => r2(28), D(27) => r2(27), D(26) 
                           => r2(26), D(25) => r2(25), D(24) => r2(24), D(23) 
                           => r2(23), D(22) => r2(22), D(21) => r2(21), D(20) 
                           => r2(20), D(19) => r2(19), D(18) => r2(18), D(17) 
                           => r2(17), D(16) => r2(16), D(15) => r2(15), D(14) 
                           => r2(14), D(13) => r2(13), D(12) => r2(12), D(11) 
                           => r2(11), D(10) => r2(10), D(9) => r2(9), D(8) => 
                           r2(8), D(7) => r2(7), D(6) => r2(6), D(5) => r2(5), 
                           D(4) => r2(4), D(3) => r2(3), D(2) => r2(2), D(1) =>
                           r2(1), D(0) => r2(0), CK => clk, Enable_n => n2, 
                           RESET_n => rst, Q(31) => r2_out(31), Q(30) => 
                           r2_out(30), Q(29) => r2_out(29), Q(28) => r2_out(28)
                           , Q(27) => r2_out(27), Q(26) => r2_out(26), Q(25) =>
                           r2_out(25), Q(24) => r2_out(24), Q(23) => r2_out(23)
                           , Q(22) => r2_out(22), Q(21) => r2_out(21), Q(20) =>
                           r2_out(20), Q(19) => r2_out(19), Q(18) => r2_out(18)
                           , Q(17) => r2_out(17), Q(16) => r2_out(16), Q(15) =>
                           r2_out(15), Q(14) => r2_out(14), Q(13) => r2_out(13)
                           , Q(12) => r2_out(12), Q(11) => r2_out(11), Q(10) =>
                           r2_out(10), Q(9) => r2_out(9), Q(8) => r2_out(8), 
                           Q(7) => r2_out(7), Q(6) => r2_out(6), Q(5) => 
                           r2_out(5), Q(4) => r2_out(4), Q(3) => r2_out(3), 
                           Q(2) => r2_out(2), Q(1) => r2_out(1), Q(0) => 
                           r2_out(0));
   pc_br : P4_ADDER_NBIT32_NBIT_PER_BLOCK4_3 port map( A(31) => imm(31), A(30) 
                           => imm(30), A(29) => imm(29), A(28) => imm(28), 
                           A(27) => imm(27), A(26) => imm(26), A(25) => imm(25)
                           , A(24) => imm(24), A(23) => imm(23), A(22) => 
                           imm(22), A(21) => imm(21), A(20) => imm(20), A(19) 
                           => imm(19), A(18) => imm(18), A(17) => imm(17), 
                           A(16) => imm(16), A(15) => imm(15), A(14) => imm(14)
                           , A(13) => imm(13), A(12) => imm(12), A(11) => 
                           imm(11), A(10) => imm(10), A(9) => imm(9), A(8) => 
                           imm(8), A(7) => imm(7), A(6) => imm(6), A(5) => 
                           imm(5), A(4) => imm(4), A(3) => imm(3), A(2) => 
                           imm(2), A(1) => imm(1), A(0) => imm(0), B(31) => 
                           pc(31), B(30) => pc(30), B(29) => pc(29), B(28) => 
                           pc(28), B(27) => pc(27), B(26) => pc(26), B(25) => 
                           pc(25), B(24) => pc(24), B(23) => pc(23), B(22) => 
                           pc(22), B(21) => pc(21), B(20) => pc(20), B(19) => 
                           pc(19), B(18) => pc(18), B(17) => pc(17), B(16) => 
                           pc(16), B(15) => pc(15), B(14) => pc(14), B(13) => 
                           pc(13), B(12) => pc(12), B(11) => pc(11), B(10) => 
                           pc(10), B(9) => pc(9), B(8) => pc(8), B(7) => pc(7),
                           B(6) => pc(6), B(5) => pc(5), B(4) => pc(4), B(3) =>
                           pc(3), B(2) => pc(2), B(1) => pc(1), B(0) => pc(0), 
                           Cin => X_Logic0_port, Cout => n_1200, Y(31) => 
                           pc_b_31_port, Y(30) => pc_b_30_port, Y(29) => 
                           pc_b_29_port, Y(28) => pc_b_28_port, Y(27) => 
                           pc_b_27_port, Y(26) => pc_b_26_port, Y(25) => 
                           pc_b_25_port, Y(24) => pc_b_24_port, Y(23) => 
                           pc_b_23_port, Y(22) => pc_b_22_port, Y(21) => 
                           pc_b_21_port, Y(20) => pc_b_20_port, Y(19) => 
                           pc_b_19_port, Y(18) => pc_b_18_port, Y(17) => 
                           pc_b_17_port, Y(16) => pc_b_16_port, Y(15) => 
                           pc_b_15_port, Y(14) => pc_b_14_port, Y(13) => 
                           pc_b_13_port, Y(12) => pc_b_12_port, Y(11) => 
                           pc_b_11_port, Y(10) => pc_b_10_port, Y(9) => 
                           pc_b_9_port, Y(8) => pc_b_8_port, Y(7) => 
                           pc_b_7_port, Y(6) => pc_b_6_port, Y(5) => 
                           pc_b_5_port, Y(4) => pc_b_4_port, Y(3) => 
                           pc_b_3_port, Y(2) => pc_b_2_port, Y(1) => 
                           pc_b_1_port, Y(0) => pc_b_0_port);
   pc_jp : P4_ADDER_NBIT32_NBIT_PER_BLOCK4_2 port map( A(31) => j_lab(31), 
                           A(30) => j_lab(30), A(29) => j_lab(29), A(28) => 
                           j_lab(28), A(27) => j_lab(27), A(26) => j_lab(26), 
                           A(25) => j_lab(25), A(24) => j_lab(24), A(23) => 
                           j_lab(23), A(22) => j_lab(22), A(21) => j_lab(21), 
                           A(20) => j_lab(20), A(19) => j_lab(19), A(18) => 
                           j_lab(18), A(17) => j_lab(17), A(16) => j_lab(16), 
                           A(15) => j_lab(15), A(14) => j_lab(14), A(13) => 
                           j_lab(13), A(12) => j_lab(12), A(11) => j_lab(11), 
                           A(10) => j_lab(10), A(9) => j_lab(9), A(8) => 
                           j_lab(8), A(7) => j_lab(7), A(6) => j_lab(6), A(5) 
                           => j_lab(5), A(4) => j_lab(4), A(3) => j_lab(3), 
                           A(2) => j_lab(2), A(1) => j_lab(1), A(0) => j_lab(0)
                           , B(31) => pc(31), B(30) => pc(30), B(29) => pc(29),
                           B(28) => pc(28), B(27) => pc(27), B(26) => pc(26), 
                           B(25) => pc(25), B(24) => pc(24), B(23) => pc(23), 
                           B(22) => pc(22), B(21) => pc(21), B(20) => pc(20), 
                           B(19) => pc(19), B(18) => pc(18), B(17) => pc(17), 
                           B(16) => pc(16), B(15) => pc(15), B(14) => pc(14), 
                           B(13) => pc(13), B(12) => pc(12), B(11) => pc(11), 
                           B(10) => pc(10), B(9) => pc(9), B(8) => pc(8), B(7) 
                           => pc(7), B(6) => pc(6), B(5) => pc(5), B(4) => 
                           pc(4), B(3) => pc(3), B(2) => pc(2), B(1) => pc(1), 
                           B(0) => pc(0), Cin => X_Logic0_port, Cout => n_1201,
                           Y(31) => pc_j_31_port, Y(30) => pc_j_30_port, Y(29) 
                           => pc_j_29_port, Y(28) => pc_j_28_port, Y(27) => 
                           pc_j_27_port, Y(26) => pc_j_26_port, Y(25) => 
                           pc_j_25_port, Y(24) => pc_j_24_port, Y(23) => 
                           pc_j_23_port, Y(22) => pc_j_22_port, Y(21) => 
                           pc_j_21_port, Y(20) => pc_j_20_port, Y(19) => 
                           pc_j_19_port, Y(18) => pc_j_18_port, Y(17) => 
                           pc_j_17_port, Y(16) => pc_j_16_port, Y(15) => 
                           pc_j_15_port, Y(14) => pc_j_14_port, Y(13) => 
                           pc_j_13_port, Y(12) => pc_j_12_port, Y(11) => 
                           pc_j_11_port, Y(10) => pc_j_10_port, Y(9) => 
                           pc_j_9_port, Y(8) => pc_j_8_port, Y(7) => 
                           pc_j_7_port, Y(6) => pc_j_6_port, Y(5) => 
                           pc_j_5_port, Y(4) => pc_j_4_port, Y(3) => 
                           pc_j_3_port, Y(2) => pc_j_2_port, Y(1) => 
                           pc_j_1_port, Y(0) => pc_j_0_port);
   pc_reg_b : REG_GEN_NBIT32_7 port map( D(31) => pc_b_31_port, D(30) => 
                           pc_b_30_port, D(29) => pc_b_29_port, D(28) => 
                           pc_b_28_port, D(27) => pc_b_27_port, D(26) => 
                           pc_b_26_port, D(25) => pc_b_25_port, D(24) => 
                           pc_b_24_port, D(23) => pc_b_23_port, D(22) => 
                           pc_b_22_port, D(21) => pc_b_21_port, D(20) => 
                           pc_b_20_port, D(19) => pc_b_19_port, D(18) => 
                           pc_b_18_port, D(17) => pc_b_17_port, D(16) => 
                           pc_b_16_port, D(15) => pc_b_15_port, D(14) => 
                           pc_b_14_port, D(13) => pc_b_13_port, D(12) => 
                           pc_b_12_port, D(11) => pc_b_11_port, D(10) => 
                           pc_b_10_port, D(9) => pc_b_9_port, D(8) => 
                           pc_b_8_port, D(7) => pc_b_7_port, D(6) => 
                           pc_b_6_port, D(5) => pc_b_5_port, D(4) => 
                           pc_b_4_port, D(3) => pc_b_3_port, D(2) => 
                           pc_b_2_port, D(1) => pc_b_1_port, D(0) => 
                           pc_b_0_port, CK => clk, Enable_n => n2, RESET_n => 
                           rst, Q(31) => b_lab_out(31), Q(30) => b_lab_out(30),
                           Q(29) => b_lab_out(29), Q(28) => b_lab_out(28), 
                           Q(27) => b_lab_out(27), Q(26) => b_lab_out(26), 
                           Q(25) => b_lab_out(25), Q(24) => b_lab_out(24), 
                           Q(23) => b_lab_out(23), Q(22) => b_lab_out(22), 
                           Q(21) => b_lab_out(21), Q(20) => b_lab_out(20), 
                           Q(19) => b_lab_out(19), Q(18) => b_lab_out(18), 
                           Q(17) => b_lab_out(17), Q(16) => b_lab_out(16), 
                           Q(15) => b_lab_out(15), Q(14) => b_lab_out(14), 
                           Q(13) => b_lab_out(13), Q(12) => b_lab_out(12), 
                           Q(11) => b_lab_out(11), Q(10) => b_lab_out(10), Q(9)
                           => b_lab_out(9), Q(8) => b_lab_out(8), Q(7) => 
                           b_lab_out(7), Q(6) => b_lab_out(6), Q(5) => 
                           b_lab_out(5), Q(4) => b_lab_out(4), Q(3) => 
                           b_lab_out(3), Q(2) => b_lab_out(2), Q(1) => 
                           b_lab_out(1), Q(0) => b_lab_out(0));
   pc_reg_j : REG_GEN_NBIT32_6 port map( D(31) => pc_j_31_port, D(30) => 
                           pc_j_30_port, D(29) => pc_j_29_port, D(28) => 
                           pc_j_28_port, D(27) => pc_j_27_port, D(26) => 
                           pc_j_26_port, D(25) => pc_j_25_port, D(24) => 
                           pc_j_24_port, D(23) => pc_j_23_port, D(22) => 
                           pc_j_22_port, D(21) => pc_j_21_port, D(20) => 
                           pc_j_20_port, D(19) => pc_j_19_port, D(18) => 
                           pc_j_18_port, D(17) => pc_j_17_port, D(16) => 
                           pc_j_16_port, D(15) => pc_j_15_port, D(14) => 
                           pc_j_14_port, D(13) => pc_j_13_port, D(12) => 
                           pc_j_12_port, D(11) => pc_j_11_port, D(10) => 
                           pc_j_10_port, D(9) => pc_j_9_port, D(8) => 
                           pc_j_8_port, D(7) => pc_j_7_port, D(6) => 
                           pc_j_6_port, D(5) => pc_j_5_port, D(4) => 
                           pc_j_4_port, D(3) => pc_j_3_port, D(2) => 
                           pc_j_2_port, D(1) => pc_j_1_port, D(0) => 
                           pc_j_0_port, CK => clk, Enable_n => n2, RESET_n => 
                           rst, Q(31) => j_lab_out(31), Q(30) => j_lab_out(30),
                           Q(29) => j_lab_out(29), Q(28) => j_lab_out(28), 
                           Q(27) => j_lab_out(27), Q(26) => j_lab_out(26), 
                           Q(25) => j_lab_out(25), Q(24) => j_lab_out(24), 
                           Q(23) => j_lab_out(23), Q(22) => j_lab_out(22), 
                           Q(21) => j_lab_out(21), Q(20) => j_lab_out(20), 
                           Q(19) => j_lab_out(19), Q(18) => j_lab_out(18), 
                           Q(17) => j_lab_out(17), Q(16) => j_lab_out(16), 
                           Q(15) => j_lab_out(15), Q(14) => j_lab_out(14), 
                           Q(13) => j_lab_out(13), Q(12) => j_lab_out(12), 
                           Q(11) => j_lab_out(11), Q(10) => j_lab_out(10), Q(9)
                           => j_lab_out(9), Q(8) => j_lab_out(8), Q(7) => 
                           j_lab_out(7), Q(6) => j_lab_out(6), Q(5) => 
                           j_lab_out(5), Q(4) => j_lab_out(4), Q(3) => 
                           j_lab_out(3), Q(2) => j_lab_out(2), Q(1) => 
                           j_lab_out(1), Q(0) => j_lab_out(0));
   pc_reg : REG_GEN_NBIT32_5 port map( D(31) => pc(31), D(30) => pc(30), D(29) 
                           => pc(29), D(28) => pc(28), D(27) => pc(27), D(26) 
                           => pc(26), D(25) => pc(25), D(24) => pc(24), D(23) 
                           => pc(23), D(22) => pc(22), D(21) => pc(21), D(20) 
                           => pc(20), D(19) => pc(19), D(18) => pc(18), D(17) 
                           => pc(17), D(16) => pc(16), D(15) => pc(15), D(14) 
                           => pc(14), D(13) => pc(13), D(12) => pc(12), D(11) 
                           => pc(11), D(10) => pc(10), D(9) => pc(9), D(8) => 
                           pc(8), D(7) => pc(7), D(6) => pc(6), D(5) => pc(5), 
                           D(4) => pc(4), D(3) => pc(3), D(2) => pc(2), D(1) =>
                           pc(1), D(0) => pc(0), CK => clk, Enable_n => n2, 
                           RESET_n => rst, Q(31) => pc_exe_out(31), Q(30) => 
                           pc_exe_out(30), Q(29) => pc_exe_out(29), Q(28) => 
                           pc_exe_out(28), Q(27) => pc_exe_out(27), Q(26) => 
                           pc_exe_out(26), Q(25) => pc_exe_out(25), Q(24) => 
                           pc_exe_out(24), Q(23) => pc_exe_out(23), Q(22) => 
                           pc_exe_out(22), Q(21) => pc_exe_out(21), Q(20) => 
                           pc_exe_out(20), Q(19) => pc_exe_out(19), Q(18) => 
                           pc_exe_out(18), Q(17) => pc_exe_out(17), Q(16) => 
                           pc_exe_out(16), Q(15) => pc_exe_out(15), Q(14) => 
                           pc_exe_out(14), Q(13) => pc_exe_out(13), Q(12) => 
                           pc_exe_out(12), Q(11) => pc_exe_out(11), Q(10) => 
                           pc_exe_out(10), Q(9) => pc_exe_out(9), Q(8) => 
                           pc_exe_out(8), Q(7) => pc_exe_out(7), Q(6) => 
                           pc_exe_out(6), Q(5) => pc_exe_out(5), Q(4) => 
                           pc_exe_out(4), Q(3) => pc_exe_out(3), Q(2) => 
                           pc_exe_out(2), Q(1) => pc_exe_out(1), Q(0) => 
                           pc_exe_out(0));
   rw_reg : REG_GEN_NBIT32_4 port map( D(31) => rw_s_31_port, D(30) => 
                           rw_s_30_port, D(29) => rw_s_29_port, D(28) => 
                           rw_s_28_port, D(27) => rw_s_27_port, D(26) => 
                           rw_s_26_port, D(25) => rw_s_25_port, D(24) => 
                           rw_s_24_port, D(23) => rw_s_23_port, D(22) => 
                           rw_s_22_port, D(21) => rw_s_21_port, D(20) => 
                           rw_s_20_port, D(19) => rw_s_19_port, D(18) => 
                           rw_s_18_port, D(17) => rw_s_17_port, D(16) => 
                           rw_s_16_port, D(15) => rw_s_15_port, D(14) => 
                           rw_s_14_port, D(13) => rw_s_13_port, D(12) => 
                           rw_s_12_port, D(11) => rw_s_11_port, D(10) => 
                           rw_s_10_port, D(9) => rw_s_9_port, D(8) => 
                           rw_s_8_port, D(7) => rw_s_7_port, D(6) => 
                           rw_s_6_port, D(5) => rw_s_5_port, D(4) => 
                           rw_s_4_port, D(3) => rw_s_3_port, D(2) => 
                           rw_s_2_port, D(1) => rw_s_1_port, D(0) => 
                           rw_s_0_port, CK => clk, Enable_n => n2, RESET_n => 
                           rst, Q(31) => rw_exe(31), Q(30) => rw_exe(30), Q(29)
                           => rw_exe(29), Q(28) => rw_exe(28), Q(27) => 
                           rw_exe(27), Q(26) => rw_exe(26), Q(25) => rw_exe(25)
                           , Q(24) => rw_exe(24), Q(23) => rw_exe(23), Q(22) =>
                           rw_exe(22), Q(21) => rw_exe(21), Q(20) => rw_exe(20)
                           , Q(19) => rw_exe(19), Q(18) => rw_exe(18), Q(17) =>
                           rw_exe(17), Q(16) => rw_exe(16), Q(15) => rw_exe(15)
                           , Q(14) => rw_exe(14), Q(13) => rw_exe(13), Q(12) =>
                           rw_exe(12), Q(11) => rw_exe(11), Q(10) => rw_exe(10)
                           , Q(9) => rw_exe(9), Q(8) => rw_exe(8), Q(7) => 
                           rw_exe(7), Q(6) => rw_exe(6), Q(5) => rw_exe(5), 
                           Q(4) => rw_exe(4), Q(3) => rw_exe(3), Q(2) => 
                           rw_exe(2), Q(1) => rw_exe(1), Q(0) => rw_exe(0));
   U2 : BUF_X1 port map( A => r1(25), Z => n1);
   U3 : BUF_X1 port map( A => en_reg, Z => n2);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity decodeUnit_nbit32 is

   port( Clk, Rst, en_reg, RD1, RD2 : in std_logic;  IRAM_instr, PC_Next : in 
         std_logic_vector (31 downto 0);  WR : in std_logic;  ADD_RW : in 
         std_logic_vector (4 downto 0);  DATA_RW : in std_logic_vector (31 
         downto 0);  RW_R_out, RW_I_out, Jump_address, I_immediate_ext_out, 
         RD_data_1_out, RD_data_2_out, PC_Next_out : out std_logic_vector (31 
         downto 0);  Opcode : out std_logic_vector (5 downto 0);  Func : out 
         std_logic_vector (10 downto 0));

end decodeUnit_nbit32;

architecture SYN_Behavioral of decodeUnit_nbit32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component REG_GEN_NBIT32_10
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_11
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_12
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_13
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_14
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_15
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_16
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_extension_sign_init16_sign_ext32
      port( data_in : in std_logic_vector (15 downto 0);  data_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component register_file_nbit_reg32_n_reg32_nbit_addr5
      port( reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, 
            add_rd2 : in std_logic_vector (4 downto 0);  datain : in 
            std_logic_vector (31 downto 0);  out1, out2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component sign_extension_sign_init26_sign_ext32
      port( data_in : in std_logic_vector (25 downto 0);  data_out : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, Jump_addr_31_port, Jump_addr_30_port, 
      Jump_addr_29_port, Jump_addr_28_port, Jump_addr_27_port, 
      Jump_addr_26_port, Jump_addr_25_port, Jump_addr_24_port, 
      Jump_addr_23_port, Jump_addr_22_port, Jump_addr_21_port, 
      Jump_addr_20_port, Jump_addr_19_port, Jump_addr_18_port, 
      Jump_addr_17_port, Jump_addr_16_port, Jump_addr_15_port, 
      Jump_addr_14_port, Jump_addr_13_port, Jump_addr_12_port, 
      Jump_addr_11_port, Jump_addr_10_port, Jump_addr_9_port, Jump_addr_8_port,
      Jump_addr_7_port, Jump_addr_6_port, Jump_addr_5_port, Jump_addr_4_port, 
      Jump_addr_3_port, Jump_addr_2_port, Jump_addr_1_port, Jump_addr_0_port, 
      RD_data_1_31_port, RD_data_1_30_port, RD_data_1_29_port, 
      RD_data_1_28_port, RD_data_1_27_port, RD_data_1_26_port, 
      RD_data_1_25_port, RD_data_1_24_port, RD_data_1_23_port, 
      RD_data_1_22_port, RD_data_1_21_port, RD_data_1_20_port, 
      RD_data_1_19_port, RD_data_1_18_port, RD_data_1_17_port, 
      RD_data_1_16_port, RD_data_1_15_port, RD_data_1_14_port, 
      RD_data_1_13_port, RD_data_1_12_port, RD_data_1_11_port, 
      RD_data_1_10_port, RD_data_1_9_port, RD_data_1_8_port, RD_data_1_7_port, 
      RD_data_1_6_port, RD_data_1_5_port, RD_data_1_4_port, RD_data_1_3_port, 
      RD_data_1_2_port, RD_data_1_1_port, RD_data_1_0_port, RD_data_2_31_port, 
      RD_data_2_30_port, RD_data_2_29_port, RD_data_2_28_port, 
      RD_data_2_27_port, RD_data_2_26_port, RD_data_2_25_port, 
      RD_data_2_24_port, RD_data_2_23_port, RD_data_2_22_port, 
      RD_data_2_21_port, RD_data_2_20_port, RD_data_2_19_port, 
      RD_data_2_18_port, RD_data_2_17_port, RD_data_2_16_port, 
      RD_data_2_15_port, RD_data_2_14_port, RD_data_2_13_port, 
      RD_data_2_12_port, RD_data_2_11_port, RD_data_2_10_port, RD_data_2_9_port
      , RD_data_2_8_port, RD_data_2_7_port, RD_data_2_6_port, RD_data_2_5_port,
      RD_data_2_4_port, RD_data_2_3_port, RD_data_2_2_port, RD_data_2_1_port, 
      RD_data_2_0_port, I_immediate_ext_31_port, I_immediate_ext_30_port, 
      I_immediate_ext_29_port, I_immediate_ext_28_port, I_immediate_ext_27_port
      , I_immediate_ext_26_port, I_immediate_ext_25_port, 
      I_immediate_ext_24_port, I_immediate_ext_23_port, I_immediate_ext_22_port
      , I_immediate_ext_21_port, I_immediate_ext_20_port, 
      I_immediate_ext_19_port, I_immediate_ext_18_port, I_immediate_ext_17_port
      , I_immediate_ext_16_port, I_immediate_ext_15_port, 
      I_immediate_ext_14_port, I_immediate_ext_13_port, I_immediate_ext_12_port
      , I_immediate_ext_11_port, I_immediate_ext_10_port, 
      I_immediate_ext_9_port, I_immediate_ext_8_port, I_immediate_ext_7_port, 
      I_immediate_ext_6_port, I_immediate_ext_5_port, I_immediate_ext_4_port, 
      I_immediate_ext_3_port, I_immediate_ext_2_port, I_immediate_ext_1_port, 
      I_immediate_ext_0_port, n1 : std_logic;

begin
   Opcode <= ( IRAM_instr(31), IRAM_instr(30), IRAM_instr(29), IRAM_instr(28), 
      IRAM_instr(27), IRAM_instr(26) );
   Func <= ( IRAM_instr(10), IRAM_instr(9), IRAM_instr(8), IRAM_instr(7), 
      IRAM_instr(6), IRAM_instr(5), IRAM_instr(4), IRAM_instr(3), IRAM_instr(2)
      , IRAM_instr(1), IRAM_instr(0) );
   
   X_Logic0_port <= '0';
   SIGN_EXT_immediate_J : sign_extension_sign_init26_sign_ext32 port map( 
                           data_in(25) => IRAM_instr(25), data_in(24) => 
                           IRAM_instr(24), data_in(23) => IRAM_instr(23), 
                           data_in(22) => IRAM_instr(22), data_in(21) => 
                           IRAM_instr(21), data_in(20) => IRAM_instr(20), 
                           data_in(19) => IRAM_instr(19), data_in(18) => 
                           IRAM_instr(18), data_in(17) => IRAM_instr(17), 
                           data_in(16) => IRAM_instr(16), data_in(15) => 
                           IRAM_instr(15), data_in(14) => IRAM_instr(14), 
                           data_in(13) => IRAM_instr(13), data_in(12) => 
                           IRAM_instr(12), data_in(11) => IRAM_instr(11), 
                           data_in(10) => IRAM_instr(10), data_in(9) => 
                           IRAM_instr(9), data_in(8) => IRAM_instr(8), 
                           data_in(7) => IRAM_instr(7), data_in(6) => 
                           IRAM_instr(6), data_in(5) => IRAM_instr(5), 
                           data_in(4) => IRAM_instr(4), data_in(3) => 
                           IRAM_instr(3), data_in(2) => IRAM_instr(2), 
                           data_in(1) => IRAM_instr(1), data_in(0) => 
                           IRAM_instr(0), data_out(31) => Jump_addr_31_port, 
                           data_out(30) => Jump_addr_30_port, data_out(29) => 
                           Jump_addr_29_port, data_out(28) => Jump_addr_28_port
                           , data_out(27) => Jump_addr_27_port, data_out(26) =>
                           Jump_addr_26_port, data_out(25) => Jump_addr_25_port
                           , data_out(24) => Jump_addr_24_port, data_out(23) =>
                           Jump_addr_23_port, data_out(22) => Jump_addr_22_port
                           , data_out(21) => Jump_addr_21_port, data_out(20) =>
                           Jump_addr_20_port, data_out(19) => Jump_addr_19_port
                           , data_out(18) => Jump_addr_18_port, data_out(17) =>
                           Jump_addr_17_port, data_out(16) => Jump_addr_16_port
                           , data_out(15) => Jump_addr_15_port, data_out(14) =>
                           Jump_addr_14_port, data_out(13) => Jump_addr_13_port
                           , data_out(12) => Jump_addr_12_port, data_out(11) =>
                           Jump_addr_11_port, data_out(10) => Jump_addr_10_port
                           , data_out(9) => Jump_addr_9_port, data_out(8) => 
                           Jump_addr_8_port, data_out(7) => Jump_addr_7_port, 
                           data_out(6) => Jump_addr_6_port, data_out(5) => 
                           Jump_addr_5_port, data_out(4) => Jump_addr_4_port, 
                           data_out(3) => Jump_addr_3_port, data_out(2) => 
                           Jump_addr_2_port, data_out(1) => Jump_addr_1_port, 
                           data_out(0) => Jump_addr_0_port);
   REGISTERS : register_file_nbit_reg32_n_reg32_nbit_addr5 port map( reset => 
                           Rst, enable => X_Logic0_port, rd1 => RD1, rd2 => RD2
                           , wr => WR, add_wr(4) => ADD_RW(4), add_wr(3) => 
                           ADD_RW(3), add_wr(2) => ADD_RW(2), add_wr(1) => 
                           ADD_RW(1), add_wr(0) => ADD_RW(0), add_rd1(4) => 
                           IRAM_instr(25), add_rd1(3) => IRAM_instr(24), 
                           add_rd1(2) => IRAM_instr(23), add_rd1(1) => 
                           IRAM_instr(22), add_rd1(0) => IRAM_instr(21), 
                           add_rd2(4) => IRAM_instr(20), add_rd2(3) => 
                           IRAM_instr(19), add_rd2(2) => IRAM_instr(18), 
                           add_rd2(1) => IRAM_instr(17), add_rd2(0) => 
                           IRAM_instr(16), datain(31) => DATA_RW(31), 
                           datain(30) => DATA_RW(30), datain(29) => DATA_RW(29)
                           , datain(28) => DATA_RW(28), datain(27) => 
                           DATA_RW(27), datain(26) => DATA_RW(26), datain(25) 
                           => DATA_RW(25), datain(24) => DATA_RW(24), 
                           datain(23) => DATA_RW(23), datain(22) => DATA_RW(22)
                           , datain(21) => DATA_RW(21), datain(20) => 
                           DATA_RW(20), datain(19) => DATA_RW(19), datain(18) 
                           => DATA_RW(18), datain(17) => DATA_RW(17), 
                           datain(16) => DATA_RW(16), datain(15) => DATA_RW(15)
                           , datain(14) => DATA_RW(14), datain(13) => 
                           DATA_RW(13), datain(12) => DATA_RW(12), datain(11) 
                           => DATA_RW(11), datain(10) => DATA_RW(10), datain(9)
                           => DATA_RW(9), datain(8) => DATA_RW(8), datain(7) =>
                           DATA_RW(7), datain(6) => DATA_RW(6), datain(5) => 
                           DATA_RW(5), datain(4) => DATA_RW(4), datain(3) => 
                           DATA_RW(3), datain(2) => DATA_RW(2), datain(1) => 
                           DATA_RW(1), datain(0) => DATA_RW(0), out1(31) => 
                           RD_data_1_31_port, out1(30) => RD_data_1_30_port, 
                           out1(29) => RD_data_1_29_port, out1(28) => 
                           RD_data_1_28_port, out1(27) => RD_data_1_27_port, 
                           out1(26) => RD_data_1_26_port, out1(25) => 
                           RD_data_1_25_port, out1(24) => RD_data_1_24_port, 
                           out1(23) => RD_data_1_23_port, out1(22) => 
                           RD_data_1_22_port, out1(21) => RD_data_1_21_port, 
                           out1(20) => RD_data_1_20_port, out1(19) => 
                           RD_data_1_19_port, out1(18) => RD_data_1_18_port, 
                           out1(17) => RD_data_1_17_port, out1(16) => 
                           RD_data_1_16_port, out1(15) => RD_data_1_15_port, 
                           out1(14) => RD_data_1_14_port, out1(13) => 
                           RD_data_1_13_port, out1(12) => RD_data_1_12_port, 
                           out1(11) => RD_data_1_11_port, out1(10) => 
                           RD_data_1_10_port, out1(9) => RD_data_1_9_port, 
                           out1(8) => RD_data_1_8_port, out1(7) => 
                           RD_data_1_7_port, out1(6) => RD_data_1_6_port, 
                           out1(5) => RD_data_1_5_port, out1(4) => 
                           RD_data_1_4_port, out1(3) => RD_data_1_3_port, 
                           out1(2) => RD_data_1_2_port, out1(1) => 
                           RD_data_1_1_port, out1(0) => RD_data_1_0_port, 
                           out2(31) => RD_data_2_31_port, out2(30) => 
                           RD_data_2_30_port, out2(29) => RD_data_2_29_port, 
                           out2(28) => RD_data_2_28_port, out2(27) => 
                           RD_data_2_27_port, out2(26) => RD_data_2_26_port, 
                           out2(25) => RD_data_2_25_port, out2(24) => 
                           RD_data_2_24_port, out2(23) => RD_data_2_23_port, 
                           out2(22) => RD_data_2_22_port, out2(21) => 
                           RD_data_2_21_port, out2(20) => RD_data_2_20_port, 
                           out2(19) => RD_data_2_19_port, out2(18) => 
                           RD_data_2_18_port, out2(17) => RD_data_2_17_port, 
                           out2(16) => RD_data_2_16_port, out2(15) => 
                           RD_data_2_15_port, out2(14) => RD_data_2_14_port, 
                           out2(13) => RD_data_2_13_port, out2(12) => 
                           RD_data_2_12_port, out2(11) => RD_data_2_11_port, 
                           out2(10) => RD_data_2_10_port, out2(9) => 
                           RD_data_2_9_port, out2(8) => RD_data_2_8_port, 
                           out2(7) => RD_data_2_7_port, out2(6) => 
                           RD_data_2_6_port, out2(5) => RD_data_2_5_port, 
                           out2(4) => RD_data_2_4_port, out2(3) => 
                           RD_data_2_3_port, out2(2) => RD_data_2_2_port, 
                           out2(1) => RD_data_2_1_port, out2(0) => 
                           RD_data_2_0_port);
   SIGN_EXT_immediate_I : sign_extension_sign_init16_sign_ext32 port map( 
                           data_in(15) => IRAM_instr(15), data_in(14) => 
                           IRAM_instr(14), data_in(13) => IRAM_instr(13), 
                           data_in(12) => IRAM_instr(12), data_in(11) => 
                           IRAM_instr(11), data_in(10) => IRAM_instr(10), 
                           data_in(9) => IRAM_instr(9), data_in(8) => 
                           IRAM_instr(8), data_in(7) => IRAM_instr(7), 
                           data_in(6) => IRAM_instr(6), data_in(5) => 
                           IRAM_instr(5), data_in(4) => IRAM_instr(4), 
                           data_in(3) => IRAM_instr(3), data_in(2) => 
                           IRAM_instr(2), data_in(1) => IRAM_instr(1), 
                           data_in(0) => IRAM_instr(0), data_out(31) => 
                           I_immediate_ext_31_port, data_out(30) => 
                           I_immediate_ext_30_port, data_out(29) => 
                           I_immediate_ext_29_port, data_out(28) => 
                           I_immediate_ext_28_port, data_out(27) => 
                           I_immediate_ext_27_port, data_out(26) => 
                           I_immediate_ext_26_port, data_out(25) => 
                           I_immediate_ext_25_port, data_out(24) => 
                           I_immediate_ext_24_port, data_out(23) => 
                           I_immediate_ext_23_port, data_out(22) => 
                           I_immediate_ext_22_port, data_out(21) => 
                           I_immediate_ext_21_port, data_out(20) => 
                           I_immediate_ext_20_port, data_out(19) => 
                           I_immediate_ext_19_port, data_out(18) => 
                           I_immediate_ext_18_port, data_out(17) => 
                           I_immediate_ext_17_port, data_out(16) => 
                           I_immediate_ext_16_port, data_out(15) => 
                           I_immediate_ext_15_port, data_out(14) => 
                           I_immediate_ext_14_port, data_out(13) => 
                           I_immediate_ext_13_port, data_out(12) => 
                           I_immediate_ext_12_port, data_out(11) => 
                           I_immediate_ext_11_port, data_out(10) => 
                           I_immediate_ext_10_port, data_out(9) => 
                           I_immediate_ext_9_port, data_out(8) => 
                           I_immediate_ext_8_port, data_out(7) => 
                           I_immediate_ext_7_port, data_out(6) => 
                           I_immediate_ext_6_port, data_out(5) => 
                           I_immediate_ext_5_port, data_out(4) => 
                           I_immediate_ext_4_port, data_out(3) => 
                           I_immediate_ext_3_port, data_out(2) => 
                           I_immediate_ext_2_port, data_out(1) => 
                           I_immediate_ext_1_port, data_out(0) => 
                           I_immediate_ext_0_port);
   ID_reg_RW_R : REG_GEN_NBIT32_16 port map( D(31) => X_Logic0_port, D(30) => 
                           X_Logic0_port, D(29) => X_Logic0_port, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           IRAM_instr(15), D(3) => IRAM_instr(14), D(2) => 
                           IRAM_instr(13), D(1) => IRAM_instr(12), D(0) => 
                           IRAM_instr(11), CK => Clk, Enable_n => n1, RESET_n 
                           => Rst, Q(31) => RW_R_out(31), Q(30) => RW_R_out(30)
                           , Q(29) => RW_R_out(29), Q(28) => RW_R_out(28), 
                           Q(27) => RW_R_out(27), Q(26) => RW_R_out(26), Q(25) 
                           => RW_R_out(25), Q(24) => RW_R_out(24), Q(23) => 
                           RW_R_out(23), Q(22) => RW_R_out(22), Q(21) => 
                           RW_R_out(21), Q(20) => RW_R_out(20), Q(19) => 
                           RW_R_out(19), Q(18) => RW_R_out(18), Q(17) => 
                           RW_R_out(17), Q(16) => RW_R_out(16), Q(15) => 
                           RW_R_out(15), Q(14) => RW_R_out(14), Q(13) => 
                           RW_R_out(13), Q(12) => RW_R_out(12), Q(11) => 
                           RW_R_out(11), Q(10) => RW_R_out(10), Q(9) => 
                           RW_R_out(9), Q(8) => RW_R_out(8), Q(7) => 
                           RW_R_out(7), Q(6) => RW_R_out(6), Q(5) => 
                           RW_R_out(5), Q(4) => RW_R_out(4), Q(3) => 
                           RW_R_out(3), Q(2) => RW_R_out(2), Q(1) => 
                           RW_R_out(1), Q(0) => RW_R_out(0));
   ID_reg_RW_I : REG_GEN_NBIT32_15 port map( D(31) => X_Logic0_port, D(30) => 
                           X_Logic0_port, D(29) => X_Logic0_port, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           IRAM_instr(20), D(3) => IRAM_instr(19), D(2) => 
                           IRAM_instr(18), D(1) => IRAM_instr(17), D(0) => 
                           IRAM_instr(16), CK => Clk, Enable_n => n1, RESET_n 
                           => Rst, Q(31) => RW_I_out(31), Q(30) => RW_I_out(30)
                           , Q(29) => RW_I_out(29), Q(28) => RW_I_out(28), 
                           Q(27) => RW_I_out(27), Q(26) => RW_I_out(26), Q(25) 
                           => RW_I_out(25), Q(24) => RW_I_out(24), Q(23) => 
                           RW_I_out(23), Q(22) => RW_I_out(22), Q(21) => 
                           RW_I_out(21), Q(20) => RW_I_out(20), Q(19) => 
                           RW_I_out(19), Q(18) => RW_I_out(18), Q(17) => 
                           RW_I_out(17), Q(16) => RW_I_out(16), Q(15) => 
                           RW_I_out(15), Q(14) => RW_I_out(14), Q(13) => 
                           RW_I_out(13), Q(12) => RW_I_out(12), Q(11) => 
                           RW_I_out(11), Q(10) => RW_I_out(10), Q(9) => 
                           RW_I_out(9), Q(8) => RW_I_out(8), Q(7) => 
                           RW_I_out(7), Q(6) => RW_I_out(6), Q(5) => 
                           RW_I_out(5), Q(4) => RW_I_out(4), Q(3) => 
                           RW_I_out(3), Q(2) => RW_I_out(2), Q(1) => 
                           RW_I_out(1), Q(0) => RW_I_out(0));
   ID_reg_I_imm : REG_GEN_NBIT32_14 port map( D(31) => I_immediate_ext_31_port,
                           D(30) => I_immediate_ext_30_port, D(29) => 
                           I_immediate_ext_29_port, D(28) => 
                           I_immediate_ext_28_port, D(27) => 
                           I_immediate_ext_27_port, D(26) => 
                           I_immediate_ext_26_port, D(25) => 
                           I_immediate_ext_25_port, D(24) => 
                           I_immediate_ext_24_port, D(23) => 
                           I_immediate_ext_23_port, D(22) => 
                           I_immediate_ext_22_port, D(21) => 
                           I_immediate_ext_21_port, D(20) => 
                           I_immediate_ext_20_port, D(19) => 
                           I_immediate_ext_19_port, D(18) => 
                           I_immediate_ext_18_port, D(17) => 
                           I_immediate_ext_17_port, D(16) => 
                           I_immediate_ext_16_port, D(15) => 
                           I_immediate_ext_15_port, D(14) => 
                           I_immediate_ext_14_port, D(13) => 
                           I_immediate_ext_13_port, D(12) => 
                           I_immediate_ext_12_port, D(11) => 
                           I_immediate_ext_11_port, D(10) => 
                           I_immediate_ext_10_port, D(9) => 
                           I_immediate_ext_9_port, D(8) => 
                           I_immediate_ext_8_port, D(7) => 
                           I_immediate_ext_7_port, D(6) => 
                           I_immediate_ext_6_port, D(5) => 
                           I_immediate_ext_5_port, D(4) => 
                           I_immediate_ext_4_port, D(3) => 
                           I_immediate_ext_3_port, D(2) => 
                           I_immediate_ext_2_port, D(1) => 
                           I_immediate_ext_1_port, D(0) => 
                           I_immediate_ext_0_port, CK => Clk, Enable_n => n1, 
                           RESET_n => Rst, Q(31) => I_immediate_ext_out(31), 
                           Q(30) => I_immediate_ext_out(30), Q(29) => 
                           I_immediate_ext_out(29), Q(28) => 
                           I_immediate_ext_out(28), Q(27) => 
                           I_immediate_ext_out(27), Q(26) => 
                           I_immediate_ext_out(26), Q(25) => 
                           I_immediate_ext_out(25), Q(24) => 
                           I_immediate_ext_out(24), Q(23) => 
                           I_immediate_ext_out(23), Q(22) => 
                           I_immediate_ext_out(22), Q(21) => 
                           I_immediate_ext_out(21), Q(20) => 
                           I_immediate_ext_out(20), Q(19) => 
                           I_immediate_ext_out(19), Q(18) => 
                           I_immediate_ext_out(18), Q(17) => 
                           I_immediate_ext_out(17), Q(16) => 
                           I_immediate_ext_out(16), Q(15) => 
                           I_immediate_ext_out(15), Q(14) => 
                           I_immediate_ext_out(14), Q(13) => 
                           I_immediate_ext_out(13), Q(12) => 
                           I_immediate_ext_out(12), Q(11) => 
                           I_immediate_ext_out(11), Q(10) => 
                           I_immediate_ext_out(10), Q(9) => 
                           I_immediate_ext_out(9), Q(8) => 
                           I_immediate_ext_out(8), Q(7) => 
                           I_immediate_ext_out(7), Q(6) => 
                           I_immediate_ext_out(6), Q(5) => 
                           I_immediate_ext_out(5), Q(4) => 
                           I_immediate_ext_out(4), Q(3) => 
                           I_immediate_ext_out(3), Q(2) => 
                           I_immediate_ext_out(2), Q(1) => 
                           I_immediate_ext_out(1), Q(0) => 
                           I_immediate_ext_out(0));
   ID_reg_J_imm : REG_GEN_NBIT32_13 port map( D(31) => Jump_addr_31_port, D(30)
                           => Jump_addr_30_port, D(29) => Jump_addr_29_port, 
                           D(28) => Jump_addr_28_port, D(27) => 
                           Jump_addr_27_port, D(26) => Jump_addr_26_port, D(25)
                           => Jump_addr_25_port, D(24) => Jump_addr_24_port, 
                           D(23) => Jump_addr_23_port, D(22) => 
                           Jump_addr_22_port, D(21) => Jump_addr_21_port, D(20)
                           => Jump_addr_20_port, D(19) => Jump_addr_19_port, 
                           D(18) => Jump_addr_18_port, D(17) => 
                           Jump_addr_17_port, D(16) => Jump_addr_16_port, D(15)
                           => Jump_addr_15_port, D(14) => Jump_addr_14_port, 
                           D(13) => Jump_addr_13_port, D(12) => 
                           Jump_addr_12_port, D(11) => Jump_addr_11_port, D(10)
                           => Jump_addr_10_port, D(9) => Jump_addr_9_port, D(8)
                           => Jump_addr_8_port, D(7) => Jump_addr_7_port, D(6) 
                           => Jump_addr_6_port, D(5) => Jump_addr_5_port, D(4) 
                           => Jump_addr_4_port, D(3) => Jump_addr_3_port, D(2) 
                           => Jump_addr_2_port, D(1) => Jump_addr_1_port, D(0) 
                           => Jump_addr_0_port, CK => Clk, Enable_n => n1, 
                           RESET_n => Rst, Q(31) => Jump_address(31), Q(30) => 
                           Jump_address(30), Q(29) => Jump_address(29), Q(28) 
                           => Jump_address(28), Q(27) => Jump_address(27), 
                           Q(26) => Jump_address(26), Q(25) => Jump_address(25)
                           , Q(24) => Jump_address(24), Q(23) => 
                           Jump_address(23), Q(22) => Jump_address(22), Q(21) 
                           => Jump_address(21), Q(20) => Jump_address(20), 
                           Q(19) => Jump_address(19), Q(18) => Jump_address(18)
                           , Q(17) => Jump_address(17), Q(16) => 
                           Jump_address(16), Q(15) => Jump_address(15), Q(14) 
                           => Jump_address(14), Q(13) => Jump_address(13), 
                           Q(12) => Jump_address(12), Q(11) => Jump_address(11)
                           , Q(10) => Jump_address(10), Q(9) => Jump_address(9)
                           , Q(8) => Jump_address(8), Q(7) => Jump_address(7), 
                           Q(6) => Jump_address(6), Q(5) => Jump_address(5), 
                           Q(4) => Jump_address(4), Q(3) => Jump_address(3), 
                           Q(2) => Jump_address(2), Q(1) => Jump_address(1), 
                           Q(0) => Jump_address(0));
   ID_reg_RD_data_1 : REG_GEN_NBIT32_12 port map( D(31) => RD_data_1_31_port, 
                           D(30) => RD_data_1_30_port, D(29) => 
                           RD_data_1_29_port, D(28) => RD_data_1_28_port, D(27)
                           => RD_data_1_27_port, D(26) => RD_data_1_26_port, 
                           D(25) => RD_data_1_25_port, D(24) => 
                           RD_data_1_24_port, D(23) => RD_data_1_23_port, D(22)
                           => RD_data_1_22_port, D(21) => RD_data_1_21_port, 
                           D(20) => RD_data_1_20_port, D(19) => 
                           RD_data_1_19_port, D(18) => RD_data_1_18_port, D(17)
                           => RD_data_1_17_port, D(16) => RD_data_1_16_port, 
                           D(15) => RD_data_1_15_port, D(14) => 
                           RD_data_1_14_port, D(13) => RD_data_1_13_port, D(12)
                           => RD_data_1_12_port, D(11) => RD_data_1_11_port, 
                           D(10) => RD_data_1_10_port, D(9) => RD_data_1_9_port
                           , D(8) => RD_data_1_8_port, D(7) => RD_data_1_7_port
                           , D(6) => RD_data_1_6_port, D(5) => RD_data_1_5_port
                           , D(4) => RD_data_1_4_port, D(3) => RD_data_1_3_port
                           , D(2) => RD_data_1_2_port, D(1) => RD_data_1_1_port
                           , D(0) => RD_data_1_0_port, CK => Clk, Enable_n => 
                           n1, RESET_n => Rst, Q(31) => RD_data_1_out(31), 
                           Q(30) => RD_data_1_out(30), Q(29) => 
                           RD_data_1_out(29), Q(28) => RD_data_1_out(28), Q(27)
                           => RD_data_1_out(27), Q(26) => RD_data_1_out(26), 
                           Q(25) => RD_data_1_out(25), Q(24) => 
                           RD_data_1_out(24), Q(23) => RD_data_1_out(23), Q(22)
                           => RD_data_1_out(22), Q(21) => RD_data_1_out(21), 
                           Q(20) => RD_data_1_out(20), Q(19) => 
                           RD_data_1_out(19), Q(18) => RD_data_1_out(18), Q(17)
                           => RD_data_1_out(17), Q(16) => RD_data_1_out(16), 
                           Q(15) => RD_data_1_out(15), Q(14) => 
                           RD_data_1_out(14), Q(13) => RD_data_1_out(13), Q(12)
                           => RD_data_1_out(12), Q(11) => RD_data_1_out(11), 
                           Q(10) => RD_data_1_out(10), Q(9) => RD_data_1_out(9)
                           , Q(8) => RD_data_1_out(8), Q(7) => RD_data_1_out(7)
                           , Q(6) => RD_data_1_out(6), Q(5) => RD_data_1_out(5)
                           , Q(4) => RD_data_1_out(4), Q(3) => RD_data_1_out(3)
                           , Q(2) => RD_data_1_out(2), Q(1) => RD_data_1_out(1)
                           , Q(0) => RD_data_1_out(0));
   ID_reg_RD_data_2 : REG_GEN_NBIT32_11 port map( D(31) => RD_data_2_31_port, 
                           D(30) => RD_data_2_30_port, D(29) => 
                           RD_data_2_29_port, D(28) => RD_data_2_28_port, D(27)
                           => RD_data_2_27_port, D(26) => RD_data_2_26_port, 
                           D(25) => RD_data_2_25_port, D(24) => 
                           RD_data_2_24_port, D(23) => RD_data_2_23_port, D(22)
                           => RD_data_2_22_port, D(21) => RD_data_2_21_port, 
                           D(20) => RD_data_2_20_port, D(19) => 
                           RD_data_2_19_port, D(18) => RD_data_2_18_port, D(17)
                           => RD_data_2_17_port, D(16) => RD_data_2_16_port, 
                           D(15) => RD_data_2_15_port, D(14) => 
                           RD_data_2_14_port, D(13) => RD_data_2_13_port, D(12)
                           => RD_data_2_12_port, D(11) => RD_data_2_11_port, 
                           D(10) => RD_data_2_10_port, D(9) => RD_data_2_9_port
                           , D(8) => RD_data_2_8_port, D(7) => RD_data_2_7_port
                           , D(6) => RD_data_2_6_port, D(5) => RD_data_2_5_port
                           , D(4) => RD_data_2_4_port, D(3) => RD_data_2_3_port
                           , D(2) => RD_data_2_2_port, D(1) => RD_data_2_1_port
                           , D(0) => RD_data_2_0_port, CK => Clk, Enable_n => 
                           n1, RESET_n => Rst, Q(31) => RD_data_2_out(31), 
                           Q(30) => RD_data_2_out(30), Q(29) => 
                           RD_data_2_out(29), Q(28) => RD_data_2_out(28), Q(27)
                           => RD_data_2_out(27), Q(26) => RD_data_2_out(26), 
                           Q(25) => RD_data_2_out(25), Q(24) => 
                           RD_data_2_out(24), Q(23) => RD_data_2_out(23), Q(22)
                           => RD_data_2_out(22), Q(21) => RD_data_2_out(21), 
                           Q(20) => RD_data_2_out(20), Q(19) => 
                           RD_data_2_out(19), Q(18) => RD_data_2_out(18), Q(17)
                           => RD_data_2_out(17), Q(16) => RD_data_2_out(16), 
                           Q(15) => RD_data_2_out(15), Q(14) => 
                           RD_data_2_out(14), Q(13) => RD_data_2_out(13), Q(12)
                           => RD_data_2_out(12), Q(11) => RD_data_2_out(11), 
                           Q(10) => RD_data_2_out(10), Q(9) => RD_data_2_out(9)
                           , Q(8) => RD_data_2_out(8), Q(7) => RD_data_2_out(7)
                           , Q(6) => RD_data_2_out(6), Q(5) => RD_data_2_out(5)
                           , Q(4) => RD_data_2_out(4), Q(3) => RD_data_2_out(3)
                           , Q(2) => RD_data_2_out(2), Q(1) => RD_data_2_out(1)
                           , Q(0) => RD_data_2_out(0));
   ID_reg_PC_next : REG_GEN_NBIT32_10 port map( D(31) => PC_Next(31), D(30) => 
                           PC_Next(30), D(29) => PC_Next(29), D(28) => 
                           PC_Next(28), D(27) => PC_Next(27), D(26) => 
                           PC_Next(26), D(25) => PC_Next(25), D(24) => 
                           PC_Next(24), D(23) => PC_Next(23), D(22) => 
                           PC_Next(22), D(21) => PC_Next(21), D(20) => 
                           PC_Next(20), D(19) => PC_Next(19), D(18) => 
                           PC_Next(18), D(17) => PC_Next(17), D(16) => 
                           PC_Next(16), D(15) => PC_Next(15), D(14) => 
                           PC_Next(14), D(13) => PC_Next(13), D(12) => 
                           PC_Next(12), D(11) => PC_Next(11), D(10) => 
                           PC_Next(10), D(9) => PC_Next(9), D(8) => PC_Next(8),
                           D(7) => PC_Next(7), D(6) => PC_Next(6), D(5) => 
                           PC_Next(5), D(4) => PC_Next(4), D(3) => PC_Next(3), 
                           D(2) => PC_Next(2), D(1) => PC_Next(1), D(0) => 
                           PC_Next(0), CK => Clk, Enable_n => n1, RESET_n => 
                           Rst, Q(31) => PC_Next_out(31), Q(30) => 
                           PC_Next_out(30), Q(29) => PC_Next_out(29), Q(28) => 
                           PC_Next_out(28), Q(27) => PC_Next_out(27), Q(26) => 
                           PC_Next_out(26), Q(25) => PC_Next_out(25), Q(24) => 
                           PC_Next_out(24), Q(23) => PC_Next_out(23), Q(22) => 
                           PC_Next_out(22), Q(21) => PC_Next_out(21), Q(20) => 
                           PC_Next_out(20), Q(19) => PC_Next_out(19), Q(18) => 
                           PC_Next_out(18), Q(17) => PC_Next_out(17), Q(16) => 
                           PC_Next_out(16), Q(15) => PC_Next_out(15), Q(14) => 
                           PC_Next_out(14), Q(13) => PC_Next_out(13), Q(12) => 
                           PC_Next_out(12), Q(11) => PC_Next_out(11), Q(10) => 
                           PC_Next_out(10), Q(9) => PC_Next_out(9), Q(8) => 
                           PC_Next_out(8), Q(7) => PC_Next_out(7), Q(6) => 
                           PC_Next_out(6), Q(5) => PC_Next_out(5), Q(4) => 
                           PC_Next_out(4), Q(3) => PC_Next_out(3), Q(2) => 
                           PC_Next_out(2), Q(1) => PC_Next_out(1), Q(0) => 
                           PC_Next_out(0));
   U2 : BUF_X1 port map( A => en_reg, Z => n1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity fetchUnit_nbit32 is

   port( Clk, Rst, en_reg : in std_logic;  PC_branch_jump, dout_IRAM : in 
         std_logic_vector (31 downto 0);  PC_op : in std_logic;  PC_Next_out, 
         addr_IRAM, IRAM_reg_out : out std_logic_vector (31 downto 0));

end fetchUnit_nbit32;

architecture SYN_Behavioral of fetchUnit_nbit32 is

   component REG_GEN_NBIT32_17
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_18
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component P4_ADDER_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic;  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component REG_GEN_NBIT32_0
      port( D : in std_logic_vector (31 downto 0);  CK, Enable_n, RESET_n : in 
            std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, addr_IRAM_31_port, addr_IRAM_30_port, 
      addr_IRAM_29_port, addr_IRAM_28_port, addr_IRAM_27_port, 
      addr_IRAM_26_port, addr_IRAM_25_port, addr_IRAM_24_port, 
      addr_IRAM_23_port, addr_IRAM_22_port, addr_IRAM_21_port, 
      addr_IRAM_20_port, addr_IRAM_19_port, addr_IRAM_18_port, 
      addr_IRAM_17_port, addr_IRAM_16_port, addr_IRAM_15_port, 
      addr_IRAM_14_port, addr_IRAM_13_port, addr_IRAM_12_port, 
      addr_IRAM_11_port, addr_IRAM_10_port, addr_IRAM_9_port, addr_IRAM_8_port,
      addr_IRAM_7_port, addr_IRAM_6_port, addr_IRAM_5_port, addr_IRAM_4_port, 
      addr_IRAM_3_port, addr_IRAM_2_port, addr_IRAM_1_port, addr_IRAM_0_port, 
      PC_Next_31_port, PC_Next_30_port, PC_Next_29_port, PC_Next_28_port, 
      PC_Next_27_port, PC_Next_26_port, PC_Next_25_port, PC_Next_24_port, 
      PC_Next_23_port, PC_Next_22_port, PC_Next_21_port, PC_Next_20_port, 
      PC_Next_19_port, PC_Next_18_port, PC_Next_17_port, PC_Next_16_port, 
      PC_Next_15_port, PC_Next_14_port, PC_Next_13_port, PC_Next_12_port, 
      PC_Next_11_port, PC_Next_10_port, PC_Next_9_port, PC_Next_8_port, 
      PC_Next_7_port, PC_Next_6_port, PC_Next_5_port, PC_Next_4_port, 
      PC_Next_3_port, PC_Next_2_port, PC_Next_1_port, PC_Next_0_port, 
      PC_in_31_port, PC_in_30_port, PC_in_29_port, PC_in_28_port, PC_in_27_port
      , PC_in_26_port, PC_in_25_port, PC_in_24_port, PC_in_23_port, 
      PC_in_22_port, PC_in_21_port, PC_in_20_port, PC_in_19_port, PC_in_18_port
      , PC_in_17_port, PC_in_16_port, PC_in_15_port, PC_in_14_port, 
      PC_in_13_port, PC_in_12_port, PC_in_11_port, PC_in_10_port, PC_in_9_port,
      PC_in_8_port, PC_in_7_port, PC_in_6_port, PC_in_5_port, PC_in_4_port, 
      PC_in_3_port, PC_in_2_port, PC_in_1_port, PC_in_0_port, n_1202 : 
      std_logic;

begin
   addr_IRAM <= ( addr_IRAM_31_port, addr_IRAM_30_port, addr_IRAM_29_port, 
      addr_IRAM_28_port, addr_IRAM_27_port, addr_IRAM_26_port, 
      addr_IRAM_25_port, addr_IRAM_24_port, addr_IRAM_23_port, 
      addr_IRAM_22_port, addr_IRAM_21_port, addr_IRAM_20_port, 
      addr_IRAM_19_port, addr_IRAM_18_port, addr_IRAM_17_port, 
      addr_IRAM_16_port, addr_IRAM_15_port, addr_IRAM_14_port, 
      addr_IRAM_13_port, addr_IRAM_12_port, addr_IRAM_11_port, 
      addr_IRAM_10_port, addr_IRAM_9_port, addr_IRAM_8_port, addr_IRAM_7_port, 
      addr_IRAM_6_port, addr_IRAM_5_port, addr_IRAM_4_port, addr_IRAM_3_port, 
      addr_IRAM_2_port, addr_IRAM_1_port, addr_IRAM_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   mux_PC : MUX21_GENERIC_NBIT32_0 port map( A(31) => PC_Next_31_port, A(30) =>
                           PC_Next_30_port, A(29) => PC_Next_29_port, A(28) => 
                           PC_Next_28_port, A(27) => PC_Next_27_port, A(26) => 
                           PC_Next_26_port, A(25) => PC_Next_25_port, A(24) => 
                           PC_Next_24_port, A(23) => PC_Next_23_port, A(22) => 
                           PC_Next_22_port, A(21) => PC_Next_21_port, A(20) => 
                           PC_Next_20_port, A(19) => PC_Next_19_port, A(18) => 
                           PC_Next_18_port, A(17) => PC_Next_17_port, A(16) => 
                           PC_Next_16_port, A(15) => PC_Next_15_port, A(14) => 
                           PC_Next_14_port, A(13) => PC_Next_13_port, A(12) => 
                           PC_Next_12_port, A(11) => PC_Next_11_port, A(10) => 
                           PC_Next_10_port, A(9) => PC_Next_9_port, A(8) => 
                           PC_Next_8_port, A(7) => PC_Next_7_port, A(6) => 
                           PC_Next_6_port, A(5) => PC_Next_5_port, A(4) => 
                           PC_Next_4_port, A(3) => PC_Next_3_port, A(2) => 
                           PC_Next_2_port, A(1) => PC_Next_1_port, A(0) => 
                           PC_Next_0_port, B(31) => PC_branch_jump(31), B(30) 
                           => PC_branch_jump(30), B(29) => PC_branch_jump(29), 
                           B(28) => PC_branch_jump(28), B(27) => 
                           PC_branch_jump(27), B(26) => PC_branch_jump(26), 
                           B(25) => PC_branch_jump(25), B(24) => 
                           PC_branch_jump(24), B(23) => PC_branch_jump(23), 
                           B(22) => PC_branch_jump(22), B(21) => 
                           PC_branch_jump(21), B(20) => PC_branch_jump(20), 
                           B(19) => PC_branch_jump(19), B(18) => 
                           PC_branch_jump(18), B(17) => PC_branch_jump(17), 
                           B(16) => PC_branch_jump(16), B(15) => 
                           PC_branch_jump(15), B(14) => PC_branch_jump(14), 
                           B(13) => PC_branch_jump(13), B(12) => 
                           PC_branch_jump(12), B(11) => PC_branch_jump(11), 
                           B(10) => PC_branch_jump(10), B(9) => 
                           PC_branch_jump(9), B(8) => PC_branch_jump(8), B(7) 
                           => PC_branch_jump(7), B(6) => PC_branch_jump(6), 
                           B(5) => PC_branch_jump(5), B(4) => PC_branch_jump(4)
                           , B(3) => PC_branch_jump(3), B(2) => 
                           PC_branch_jump(2), B(1) => PC_branch_jump(1), B(0) 
                           => PC_branch_jump(0), SEL => PC_op, Y(31) => 
                           PC_in_31_port, Y(30) => PC_in_30_port, Y(29) => 
                           PC_in_29_port, Y(28) => PC_in_28_port, Y(27) => 
                           PC_in_27_port, Y(26) => PC_in_26_port, Y(25) => 
                           PC_in_25_port, Y(24) => PC_in_24_port, Y(23) => 
                           PC_in_23_port, Y(22) => PC_in_22_port, Y(21) => 
                           PC_in_21_port, Y(20) => PC_in_20_port, Y(19) => 
                           PC_in_19_port, Y(18) => PC_in_18_port, Y(17) => 
                           PC_in_17_port, Y(16) => PC_in_16_port, Y(15) => 
                           PC_in_15_port, Y(14) => PC_in_14_port, Y(13) => 
                           PC_in_13_port, Y(12) => PC_in_12_port, Y(11) => 
                           PC_in_11_port, Y(10) => PC_in_10_port, Y(9) => 
                           PC_in_9_port, Y(8) => PC_in_8_port, Y(7) => 
                           PC_in_7_port, Y(6) => PC_in_6_port, Y(5) => 
                           PC_in_5_port, Y(4) => PC_in_4_port, Y(3) => 
                           PC_in_3_port, Y(2) => PC_in_2_port, Y(1) => 
                           PC_in_1_port, Y(0) => PC_in_0_port);
   PC_block : REG_GEN_NBIT32_0 port map( D(31) => PC_in_31_port, D(30) => 
                           PC_in_30_port, D(29) => PC_in_29_port, D(28) => 
                           PC_in_28_port, D(27) => PC_in_27_port, D(26) => 
                           PC_in_26_port, D(25) => PC_in_25_port, D(24) => 
                           PC_in_24_port, D(23) => PC_in_23_port, D(22) => 
                           PC_in_22_port, D(21) => PC_in_21_port, D(20) => 
                           PC_in_20_port, D(19) => PC_in_19_port, D(18) => 
                           PC_in_18_port, D(17) => PC_in_17_port, D(16) => 
                           PC_in_16_port, D(15) => PC_in_15_port, D(14) => 
                           PC_in_14_port, D(13) => PC_in_13_port, D(12) => 
                           PC_in_12_port, D(11) => PC_in_11_port, D(10) => 
                           PC_in_10_port, D(9) => PC_in_9_port, D(8) => 
                           PC_in_8_port, D(7) => PC_in_7_port, D(6) => 
                           PC_in_6_port, D(5) => PC_in_5_port, D(4) => 
                           PC_in_4_port, D(3) => PC_in_3_port, D(2) => 
                           PC_in_2_port, D(1) => PC_in_1_port, D(0) => 
                           PC_in_0_port, CK => Clk, Enable_n => en_reg, RESET_n
                           => Rst, Q(31) => addr_IRAM_31_port, Q(30) => 
                           addr_IRAM_30_port, Q(29) => addr_IRAM_29_port, Q(28)
                           => addr_IRAM_28_port, Q(27) => addr_IRAM_27_port, 
                           Q(26) => addr_IRAM_26_port, Q(25) => 
                           addr_IRAM_25_port, Q(24) => addr_IRAM_24_port, Q(23)
                           => addr_IRAM_23_port, Q(22) => addr_IRAM_22_port, 
                           Q(21) => addr_IRAM_21_port, Q(20) => 
                           addr_IRAM_20_port, Q(19) => addr_IRAM_19_port, Q(18)
                           => addr_IRAM_18_port, Q(17) => addr_IRAM_17_port, 
                           Q(16) => addr_IRAM_16_port, Q(15) => 
                           addr_IRAM_15_port, Q(14) => addr_IRAM_14_port, Q(13)
                           => addr_IRAM_13_port, Q(12) => addr_IRAM_12_port, 
                           Q(11) => addr_IRAM_11_port, Q(10) => 
                           addr_IRAM_10_port, Q(9) => addr_IRAM_9_port, Q(8) =>
                           addr_IRAM_8_port, Q(7) => addr_IRAM_7_port, Q(6) => 
                           addr_IRAM_6_port, Q(5) => addr_IRAM_5_port, Q(4) => 
                           addr_IRAM_4_port, Q(3) => addr_IRAM_3_port, Q(2) => 
                           addr_IRAM_2_port, Q(1) => addr_IRAM_1_port, Q(0) => 
                           addr_IRAM_0_port);
   PC_ADD : P4_ADDER_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => 
                           addr_IRAM_31_port, A(30) => addr_IRAM_30_port, A(29)
                           => addr_IRAM_29_port, A(28) => addr_IRAM_28_port, 
                           A(27) => addr_IRAM_27_port, A(26) => 
                           addr_IRAM_26_port, A(25) => addr_IRAM_25_port, A(24)
                           => addr_IRAM_24_port, A(23) => addr_IRAM_23_port, 
                           A(22) => addr_IRAM_22_port, A(21) => 
                           addr_IRAM_21_port, A(20) => addr_IRAM_20_port, A(19)
                           => addr_IRAM_19_port, A(18) => addr_IRAM_18_port, 
                           A(17) => addr_IRAM_17_port, A(16) => 
                           addr_IRAM_16_port, A(15) => addr_IRAM_15_port, A(14)
                           => addr_IRAM_14_port, A(13) => addr_IRAM_13_port, 
                           A(12) => addr_IRAM_12_port, A(11) => 
                           addr_IRAM_11_port, A(10) => addr_IRAM_10_port, A(9) 
                           => addr_IRAM_9_port, A(8) => addr_IRAM_8_port, A(7) 
                           => addr_IRAM_7_port, A(6) => addr_IRAM_6_port, A(5) 
                           => addr_IRAM_5_port, A(4) => addr_IRAM_4_port, A(3) 
                           => addr_IRAM_3_port, A(2) => addr_IRAM_2_port, A(1) 
                           => addr_IRAM_1_port, A(0) => addr_IRAM_0_port, B(31)
                           => X_Logic0_port, B(30) => X_Logic0_port, B(29) => 
                           X_Logic0_port, B(28) => X_Logic0_port, B(27) => 
                           X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
                           X_Logic0_port, B(24) => X_Logic0_port, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic1_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, Cin => 
                           X_Logic0_port, Cout => n_1202, Y(31) => 
                           PC_Next_31_port, Y(30) => PC_Next_30_port, Y(29) => 
                           PC_Next_29_port, Y(28) => PC_Next_28_port, Y(27) => 
                           PC_Next_27_port, Y(26) => PC_Next_26_port, Y(25) => 
                           PC_Next_25_port, Y(24) => PC_Next_24_port, Y(23) => 
                           PC_Next_23_port, Y(22) => PC_Next_22_port, Y(21) => 
                           PC_Next_21_port, Y(20) => PC_Next_20_port, Y(19) => 
                           PC_Next_19_port, Y(18) => PC_Next_18_port, Y(17) => 
                           PC_Next_17_port, Y(16) => PC_Next_16_port, Y(15) => 
                           PC_Next_15_port, Y(14) => PC_Next_14_port, Y(13) => 
                           PC_Next_13_port, Y(12) => PC_Next_12_port, Y(11) => 
                           PC_Next_11_port, Y(10) => PC_Next_10_port, Y(9) => 
                           PC_Next_9_port, Y(8) => PC_Next_8_port, Y(7) => 
                           PC_Next_7_port, Y(6) => PC_Next_6_port, Y(5) => 
                           PC_Next_5_port, Y(4) => PC_Next_4_port, Y(3) => 
                           PC_Next_3_port, Y(2) => PC_Next_2_port, Y(1) => 
                           PC_Next_1_port, Y(0) => PC_Next_0_port);
   IF_reg_PC_Next : REG_GEN_NBIT32_18 port map( D(31) => PC_Next_31_port, D(30)
                           => PC_Next_30_port, D(29) => PC_Next_29_port, D(28) 
                           => PC_Next_28_port, D(27) => PC_Next_27_port, D(26) 
                           => PC_Next_26_port, D(25) => PC_Next_25_port, D(24) 
                           => PC_Next_24_port, D(23) => PC_Next_23_port, D(22) 
                           => PC_Next_22_port, D(21) => PC_Next_21_port, D(20) 
                           => PC_Next_20_port, D(19) => PC_Next_19_port, D(18) 
                           => PC_Next_18_port, D(17) => PC_Next_17_port, D(16) 
                           => PC_Next_16_port, D(15) => PC_Next_15_port, D(14) 
                           => PC_Next_14_port, D(13) => PC_Next_13_port, D(12) 
                           => PC_Next_12_port, D(11) => PC_Next_11_port, D(10) 
                           => PC_Next_10_port, D(9) => PC_Next_9_port, D(8) => 
                           PC_Next_8_port, D(7) => PC_Next_7_port, D(6) => 
                           PC_Next_6_port, D(5) => PC_Next_5_port, D(4) => 
                           PC_Next_4_port, D(3) => PC_Next_3_port, D(2) => 
                           PC_Next_2_port, D(1) => PC_Next_1_port, D(0) => 
                           PC_Next_0_port, CK => Clk, Enable_n => en_reg, 
                           RESET_n => Rst, Q(31) => PC_Next_out(31), Q(30) => 
                           PC_Next_out(30), Q(29) => PC_Next_out(29), Q(28) => 
                           PC_Next_out(28), Q(27) => PC_Next_out(27), Q(26) => 
                           PC_Next_out(26), Q(25) => PC_Next_out(25), Q(24) => 
                           PC_Next_out(24), Q(23) => PC_Next_out(23), Q(22) => 
                           PC_Next_out(22), Q(21) => PC_Next_out(21), Q(20) => 
                           PC_Next_out(20), Q(19) => PC_Next_out(19), Q(18) => 
                           PC_Next_out(18), Q(17) => PC_Next_out(17), Q(16) => 
                           PC_Next_out(16), Q(15) => PC_Next_out(15), Q(14) => 
                           PC_Next_out(14), Q(13) => PC_Next_out(13), Q(12) => 
                           PC_Next_out(12), Q(11) => PC_Next_out(11), Q(10) => 
                           PC_Next_out(10), Q(9) => PC_Next_out(9), Q(8) => 
                           PC_Next_out(8), Q(7) => PC_Next_out(7), Q(6) => 
                           PC_Next_out(6), Q(5) => PC_Next_out(5), Q(4) => 
                           PC_Next_out(4), Q(3) => PC_Next_out(3), Q(2) => 
                           PC_Next_out(2), Q(1) => PC_Next_out(1), Q(0) => 
                           PC_Next_out(0));
   IF_reg_IRAM_out : REG_GEN_NBIT32_17 port map( D(31) => dout_IRAM(31), D(30) 
                           => dout_IRAM(30), D(29) => dout_IRAM(29), D(28) => 
                           dout_IRAM(28), D(27) => dout_IRAM(27), D(26) => 
                           dout_IRAM(26), D(25) => dout_IRAM(25), D(24) => 
                           dout_IRAM(24), D(23) => dout_IRAM(23), D(22) => 
                           dout_IRAM(22), D(21) => dout_IRAM(21), D(20) => 
                           dout_IRAM(20), D(19) => dout_IRAM(19), D(18) => 
                           dout_IRAM(18), D(17) => dout_IRAM(17), D(16) => 
                           dout_IRAM(16), D(15) => dout_IRAM(15), D(14) => 
                           dout_IRAM(14), D(13) => dout_IRAM(13), D(12) => 
                           dout_IRAM(12), D(11) => dout_IRAM(11), D(10) => 
                           dout_IRAM(10), D(9) => dout_IRAM(9), D(8) => 
                           dout_IRAM(8), D(7) => dout_IRAM(7), D(6) => 
                           dout_IRAM(6), D(5) => dout_IRAM(5), D(4) => 
                           dout_IRAM(4), D(3) => dout_IRAM(3), D(2) => 
                           dout_IRAM(2), D(1) => dout_IRAM(1), D(0) => 
                           dout_IRAM(0), CK => Clk, Enable_n => en_reg, RESET_n
                           => Rst, Q(31) => IRAM_reg_out(31), Q(30) => 
                           IRAM_reg_out(30), Q(29) => IRAM_reg_out(29), Q(28) 
                           => IRAM_reg_out(28), Q(27) => IRAM_reg_out(27), 
                           Q(26) => IRAM_reg_out(26), Q(25) => IRAM_reg_out(25)
                           , Q(24) => IRAM_reg_out(24), Q(23) => 
                           IRAM_reg_out(23), Q(22) => IRAM_reg_out(22), Q(21) 
                           => IRAM_reg_out(21), Q(20) => IRAM_reg_out(20), 
                           Q(19) => IRAM_reg_out(19), Q(18) => IRAM_reg_out(18)
                           , Q(17) => IRAM_reg_out(17), Q(16) => 
                           IRAM_reg_out(16), Q(15) => IRAM_reg_out(15), Q(14) 
                           => IRAM_reg_out(14), Q(13) => IRAM_reg_out(13), 
                           Q(12) => IRAM_reg_out(12), Q(11) => IRAM_reg_out(11)
                           , Q(10) => IRAM_reg_out(10), Q(9) => IRAM_reg_out(9)
                           , Q(8) => IRAM_reg_out(8), Q(7) => IRAM_reg_out(7), 
                           Q(6) => IRAM_reg_out(6), Q(5) => IRAM_reg_out(5), 
                           Q(4) => IRAM_reg_out(4), Q(3) => IRAM_reg_out(3), 
                           Q(2) => IRAM_reg_out(2), Q(1) => IRAM_reg_out(1), 
                           Q(0) => IRAM_reg_out(0));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE45_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   port( Clk, Rst, En : in std_logic;  IR_opcode : in std_logic_vector (5 
         downto 0);  IR_func : in std_logic_vector (10 downto 0);  PC_OP, 
         EN_REG_IF, EN_REG_ID, RD1, RD2, SEL_EX, EN_REG_EX, SEL_MUX_RW : out 
         std_logic;  ALU_OPCODE : out std_logic_vector (3 downto 0);  
         EN_REG_MEM, MEM_EN_MEM, RD_MEM, WR_MEM, B_OP_MEM, J_OP_MEM, JAL_OP_MEM
         , MEM_TO_REG_WB, WR : out std_logic);

end dlx_cu_MICROCODE_MEM_SIZE45_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE45_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ALU_OPCODE_3_port, ALU_OPCODE_2_port, 
      ALU_OPCODE_1_port, ALU_OPCODE_0_port, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n66, n68, n76, n80, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n65, n67
      , n69, n70, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212 : std_logic;

begin
   ALU_OPCODE <= ( ALU_OPCODE_3_port, ALU_OPCODE_2_port, ALU_OPCODE_1_port, 
      ALU_OPCODE_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   aluOpcode_3_reg_3_inst : DFFR_X1 port map( D => n68, CK => Clk, RN => n84, Q
                           => ALU_OPCODE_3_port, QN => n56);
   aluOpcode_3_reg_2_inst : DFFR_X1 port map( D => n87, CK => Clk, RN => n84, Q
                           => ALU_OPCODE_2_port, QN => n_1203);
   aluOpcode_3_reg_1_inst : DFFR_X1 port map( D => n66, CK => Clk, RN => n84, Q
                           => ALU_OPCODE_1_port, QN => n_1204);
   aluOpcode_3_reg_0_inst : DFFR_X1 port map( D => n80, CK => Clk, RN => n84, Q
                           => ALU_OPCODE_0_port, QN => n76);
   EN_REG_IF_reg : DFFS_X1 port map( D => X_Logic0_port, CK => Clk, SN => n85, 
                           Q => EN_REG_IF, QN => n_1205);
   EN_REG_ID_reg : DFFS_X1 port map( D => X_Logic0_port, CK => Clk, SN => n84, 
                           Q => EN_REG_ID, QN => n_1206);
   RD1_reg : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN => n84, Q => 
                           RD1, QN => n_1207);
   RD2_reg : DFFR_X1 port map( D => X_Logic1_port, CK => Clk, RN => n84, Q => 
                           RD2, QN => n_1208);
   cw3_reg_10_inst : DFFS_X1 port map( D => n64, CK => Clk, SN => n84, Q => 
                           EN_REG_EX, QN => n55);
   cw3_reg_9_inst : DFFS_X1 port map( D => n63, CK => Clk, SN => n84, Q => 
                           n_1209, QN => n53);
   cw3_reg_2_inst : DFFS_X1 port map( D => n62, CK => Clk, SN => n85, Q => 
                           n_1210, QN => n65);
   cw3_reg_1_inst : DFFS_X1 port map( D => n61, CK => Clk, SN => n84, Q => 
                           n_1211, QN => n67);
   cw4_reg_9_inst : DFFS_X1 port map( D => n60, CK => Clk, SN => n84, Q => 
                           MEM_EN_MEM, QN => n54);
   cw4_reg_1_inst : DFFS_X1 port map( D => n58, CK => Clk, SN => n84, Q => 
                           n_1212, QN => n69);
   WR <= '0';
   PC_OP <= '0';
   JAL_OP_MEM <= '0';
   J_OP_MEM <= '0';
   B_OP_MEM <= '0';
   WR_MEM <= '0';
   RD_MEM <= '0';
   SEL_MUX_RW <= '0';
   SEL_EX <= '0';
   U57 : OAI33_X1 port map( A1 => n24, A2 => IR_opcode(1), A3 => n25, B1 => n26
                           , B2 => n96, B3 => n94, ZN => n23);
   U58 : XOR2_X1 port map( A => n98, B => IR_opcode(4), Z => n25);
   U59 : OAI33_X1 port map( A1 => n88, A2 => IR_func(0), A3 => n29, B1 => n24, 
                           B2 => IR_opcode(0), B3 => n38, ZN => n37);
   U60 : OAI33_X1 port map( A1 => n34, A2 => IR_func(2), A3 => n103, B1 => n41,
                           B2 => IR_opcode(2), B3 => n98, ZN => n46);
   U61 : NAND3_X1 port map( A1 => n29, A2 => n47, A3 => IR_func(3), ZN => n34);
   U71 : NAND3_X1 port map( A1 => n89, A2 => n100, A3 => n47, ZN => n33);
   U72 : NAND3_X1 port map( A1 => n97, A2 => n93, A3 => n86, ZN => n39);
   U73 : NAND3_X1 port map( A1 => n86, A2 => IR_opcode(4), A3 => n52, ZN => n43
                           );
   U74 : NAND3_X1 port map( A1 => n89, A2 => n92, A3 => IR_opcode(2), ZN => n24
                           );
   cw5_reg_1_inst : DFFS_X1 port map( D => n57, CK => Clk, SN => n85, Q => 
                           MEM_TO_REG_WB, QN => n70);
   cw4_reg_2_inst : DFFS_X1 port map( D => n59, CK => Clk, SN => Rst, Q => 
                           EN_REG_MEM, QN => n83);
   U3 : INV_X1 port map( A => n28, ZN => n88);
   U4 : BUF_X1 port map( A => Rst, Z => n84);
   U5 : BUF_X1 port map( A => Rst, Z => n85);
   U6 : NOR2_X1 port map( A1 => n101, A2 => n33, ZN => n28);
   U7 : INV_X1 port map( A => n24, ZN => n86);
   U8 : INV_X1 port map( A => n34, ZN => n91);
   U9 : INV_X1 port map( A => n40, ZN => n96);
   U10 : AND2_X1 port map( A1 => n28, A2 => n29, ZN => n22);
   U11 : INV_X1 port map( A => IR_func(0), ZN => n103);
   U12 : INV_X1 port map( A => n27, ZN => n94);
   U13 : NAND2_X1 port map( A1 => n89, A2 => n92, ZN => n26);
   U14 : INV_X1 port map( A => En, ZN => n89);
   U15 : NOR4_X1 port map( A1 => IR_func(10), A2 => n96, A3 => n49, A4 => n50, 
                           ZN => n47);
   U16 : OR3_X1 port map( A1 => IR_func(7), A2 => IR_func(6), A3 => IR_func(4),
                           ZN => n49);
   U17 : NAND4_X1 port map( A1 => n93, A2 => n92, A3 => n95, A4 => n51, ZN => 
                           n50);
   U18 : NOR3_X1 port map( A1 => IR_func(8), A2 => IR_opcode(1), A3 => 
                           IR_func(9), ZN => n51);
   U19 : NOR4_X1 port map( A1 => IR_func(2), A2 => n99, A3 => n33, A4 => n102, 
                           ZN => n32);
   U20 : OAI222_X1 port map( A1 => En, A2 => n90, B1 => IR_opcode(3), B2 => n39
                           , C1 => n56, C2 => n89, ZN => n68);
   U21 : INV_X1 port map( A => n36, ZN => n90);
   U22 : NOR3_X1 port map( A1 => n97, A2 => IR_opcode(4), A3 => n95, ZN => n27)
                           ;
   U23 : OAI22_X1 port map( A1 => n40, A2 => n41, B1 => n42, B2 => n34, ZN => 
                           n36);
   U24 : NOR2_X1 port map( A1 => IR_func(0), A2 => IR_func(2), ZN => n42);
   U25 : INV_X1 port map( A => IR_func(3), ZN => n100);
   U26 : NOR2_X1 port map( A1 => n99, A2 => IR_func(1), ZN => n29);
   U27 : OAI221_X1 port map( B1 => IR_func(0), B2 => n20, C1 => n76, C2 => n89,
                           A => n21, ZN => n80);
   U28 : AOI221_X1 port map( B1 => n30, B2 => n91, C1 => n31, C2 => n28, A => 
                           n32, ZN => n20);
   U29 : AOI21_X1 port map( B1 => n22, B2 => IR_func(0), A => n23, ZN => n21);
   U30 : NOR2_X1 port map( A1 => IR_func(5), A2 => IR_func(1), ZN => n31);
   U31 : NOR2_X1 port map( A1 => IR_opcode(2), A2 => IR_opcode(0), ZN => n40);
   U32 : NAND4_X1 port map( A1 => n43, A2 => n39, A3 => n44, A4 => n45, ZN => 
                           n66);
   U33 : AOI22_X1 port map( A1 => n46, A2 => n89, B1 => En, B2 => 
                           ALU_OPCODE_1_port, ZN => n45);
   U34 : OAI21_X1 port map( B1 => n48, B2 => n29, A => n28, ZN => n44);
   U35 : INV_X1 port map( A => IR_opcode(5), ZN => n92);
   U36 : INV_X1 port map( A => IR_opcode(1), ZN => n97);
   U37 : INV_X1 port map( A => IR_opcode(3), ZN => n95);
   U38 : INV_X1 port map( A => IR_func(2), ZN => n101);
   U39 : INV_X1 port map( A => IR_func(5), ZN => n99);
   U40 : INV_X1 port map( A => IR_opcode(4), ZN => n93);
   U41 : INV_X1 port map( A => n35, ZN => n87);
   U42 : AOI221_X1 port map( B1 => n36, B2 => n89, C1 => En, C2 => 
                           ALU_OPCODE_2_port, A => n37, ZN => n35);
   U43 : AOI21_X1 port map( B1 => IR_opcode(4), B2 => n95, A => n27, ZN => n38)
                           ;
   U44 : NOR3_X1 port map( A1 => n102, A2 => IR_func(5), A3 => IR_func(0), ZN 
                           => n48);
   U45 : OAI22_X1 port map( A1 => n69, A2 => n89, B1 => n67, B2 => En, ZN => 
                           n58);
   U46 : OAI22_X1 port map( A1 => n89, A2 => n83, B1 => n65, B2 => En, ZN => 
                           n59);
   U47 : OAI22_X1 port map( A1 => n54, A2 => n89, B1 => n53, B2 => En, ZN => 
                           n60);
   U48 : OAI22_X1 port map( A1 => n70, A2 => n89, B1 => n69, B2 => En, ZN => 
                           n57);
   U49 : NAND4_X1 port map( A1 => IR_opcode(4), A2 => IR_opcode(3), A3 => n97, 
                           A4 => n92, ZN => n41);
   U50 : NOR3_X1 port map( A1 => n97, A2 => IR_opcode(3), A3 => IR_opcode(0), 
                           ZN => n52);
   U51 : NOR2_X1 port map( A1 => En, A2 => n101, ZN => n30);
   U52 : NOR2_X1 port map( A1 => n67, A2 => n89, ZN => n61);
   U53 : NOR2_X1 port map( A1 => n65, A2 => n89, ZN => n62);
   U54 : NOR2_X1 port map( A1 => n53, A2 => n89, ZN => n63);
   U55 : NOR2_X1 port map( A1 => n55, A2 => n89, ZN => n64);
   U56 : INV_X1 port map( A => IR_func(1), ZN => n102);
   U75 : INV_X1 port map( A => IR_opcode(0), ZN => n98);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity flip_flop_1 is

   port( D, CK, Enable_n, RESET_n : in std_logic;  Q : out std_logic);

end flip_flop_1;

architecture SYN_FF_ASYNCH of flip_flop_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n5 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => RESET_n, Q => Q, QN => n5
                           );
   U2 : OAI22_X1 port map( A1 => n5, A2 => n3, B1 => Enable_n, B2 => n2, ZN => 
                           n1);
   U3 : INV_X1 port map( A => Enable_n, ZN => n3);
   U4 : INV_X1 port map( A => D, ZN => n2);

end SYN_FF_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity flip_flop_0 is

   port( D, CK, Enable_n, RESET_n : in std_logic;  Q : out std_logic);

end flip_flop_0;

architecture SYN_FF_ASYNCH of flip_flop_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n4, n2, n3 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => RESET_n, Q => Q, QN => n4
                           );
   U2 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => Enable_n, B2 => n2, ZN => 
                           n1);
   U3 : INV_X1 port map( A => Enable_n, ZN => n3);
   U4 : INV_X1 port map( A => D, ZN => n2);

end SYN_FF_ASYNCH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity datapath_nbit32 is

   port( Clk, Rst, PC_op, en_reg_if, RD1, RD2 : in std_logic;  dout_IRAM : in 
         std_logic_vector (31 downto 0);  addr_IRAM : out std_logic_vector (31 
         downto 0);  en_reg_id, WR : in std_logic;  Opcode : out 
         std_logic_vector (5 downto 0);  Func : out std_logic_vector (10 downto
         0);  sel_ex, sel_mux_rw, en_reg_ex : in std_logic;  alu_sel : in 
         std_logic_vector (3 downto 0);  en_reg_mem : in std_logic;  
         dataout_from_mem : in std_logic_vector (31 downto 0);  addr_mem, 
         datain_mem : out std_logic_vector (31 downto 0);  b_op_mem, j_op_mem, 
         jal_op_mem, MemtoReg_wb : in std_logic;  pipe_out : out 
         std_logic_vector (31 downto 0));

end datapath_nbit32;

architecture SYN_Behavioral of datapath_nbit32 is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component writeBackUnit_nbit32
      port( MemtoReg : in std_logic;  ReadData, AluResult : in std_logic_vector
            (31 downto 0);  WriteData : out std_logic_vector (31 downto 0));
   end component;
   
   component memoryUnit_nbit32
      port( rst, clk, en_reg, b_op, j_op, jal_op : in std_logic;  alu_out, 
            r2_out, PC, lab_b, lab_j, rw_exe, dataout_from_mem : in 
            std_logic_vector (31 downto 0);  addr_mem, datain_mem, next_PC, 
            alu_out_mem, rw_mem, data_out : out std_logic_vector (31 downto 0)
            );
   end component;
   
   component executionUnit_nbit32
      port( r1, r2, imm, j_lab, pc, RW_R, RW_I : in std_logic_vector (31 downto
            0);  s2, s3, rst, clk, en_reg : in std_logic;  alu_sel : in 
            std_logic_vector (3 downto 0);  alu_out, alu_fw_out, r2_out, 
            b_lab_out, pc_exe_out, rw_exe, j_lab_out : out std_logic_vector (31
            downto 0));
   end component;
   
   component decodeUnit_nbit32
      port( Clk, Rst, en_reg, RD1, RD2 : in std_logic;  IRAM_instr, PC_Next : 
            in std_logic_vector (31 downto 0);  WR : in std_logic;  ADD_RW : in
            std_logic_vector (4 downto 0);  DATA_RW : in std_logic_vector (31 
            downto 0);  RW_R_out, RW_I_out, Jump_address, I_immediate_ext_out, 
            RD_data_1_out, RD_data_2_out, PC_Next_out : out std_logic_vector 
            (31 downto 0);  Opcode : out std_logic_vector (5 downto 0);  Func :
            out std_logic_vector (10 downto 0));
   end component;
   
   component fetchUnit_nbit32
      port( Clk, Rst, en_reg : in std_logic;  PC_branch_jump, dout_IRAM : in 
            std_logic_vector (31 downto 0);  PC_op : in std_logic;  PC_Next_out
            , addr_IRAM, IRAM_reg_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal pipe_out_31_port, pipe_out_30_port, pipe_out_29_port, 
      pipe_out_28_port, pipe_out_27_port, pipe_out_26_port, pipe_out_25_port, 
      pipe_out_24_port, pipe_out_23_port, pipe_out_22_port, pipe_out_21_port, 
      pipe_out_20_port, pipe_out_19_port, pipe_out_18_port, pipe_out_17_port, 
      pipe_out_16_port, pipe_out_15_port, pipe_out_14_port, pipe_out_13_port, 
      pipe_out_12_port, pipe_out_11_port, pipe_out_10_port, pipe_out_9_port, 
      pipe_out_8_port, pipe_out_7_port, pipe_out_6_port, pipe_out_5_port, 
      pipe_out_4_port, pipe_out_3_port, pipe_out_2_port, pipe_out_1_port, 
      pipe_out_0_port, pc_from_mem_to_fetch_31_port, 
      pc_from_mem_to_fetch_30_port, pc_from_mem_to_fetch_29_port, 
      pc_from_mem_to_fetch_28_port, pc_from_mem_to_fetch_27_port, 
      pc_from_mem_to_fetch_26_port, pc_from_mem_to_fetch_25_port, 
      pc_from_mem_to_fetch_24_port, pc_from_mem_to_fetch_23_port, 
      pc_from_mem_to_fetch_22_port, pc_from_mem_to_fetch_21_port, 
      pc_from_mem_to_fetch_20_port, pc_from_mem_to_fetch_19_port, 
      pc_from_mem_to_fetch_18_port, pc_from_mem_to_fetch_17_port, 
      pc_from_mem_to_fetch_16_port, pc_from_mem_to_fetch_15_port, 
      pc_from_mem_to_fetch_14_port, pc_from_mem_to_fetch_13_port, 
      pc_from_mem_to_fetch_12_port, pc_from_mem_to_fetch_11_port, 
      pc_from_mem_to_fetch_10_port, pc_from_mem_to_fetch_9_port, 
      pc_from_mem_to_fetch_8_port, pc_from_mem_to_fetch_7_port, 
      pc_from_mem_to_fetch_6_port, pc_from_mem_to_fetch_5_port, 
      pc_from_mem_to_fetch_4_port, pc_from_mem_to_fetch_3_port, 
      pc_from_mem_to_fetch_2_port, pc_from_mem_to_fetch_1_port, 
      pc_from_mem_to_fetch_0_port, PC_Next_fetch_31_port, PC_Next_fetch_30_port
      , PC_Next_fetch_29_port, PC_Next_fetch_28_port, PC_Next_fetch_27_port, 
      PC_Next_fetch_26_port, PC_Next_fetch_25_port, PC_Next_fetch_24_port, 
      PC_Next_fetch_23_port, PC_Next_fetch_22_port, PC_Next_fetch_21_port, 
      PC_Next_fetch_20_port, PC_Next_fetch_19_port, PC_Next_fetch_18_port, 
      PC_Next_fetch_17_port, PC_Next_fetch_16_port, PC_Next_fetch_15_port, 
      PC_Next_fetch_14_port, PC_Next_fetch_13_port, PC_Next_fetch_12_port, 
      PC_Next_fetch_11_port, PC_Next_fetch_10_port, PC_Next_fetch_9_port, 
      PC_Next_fetch_8_port, PC_Next_fetch_7_port, PC_Next_fetch_6_port, 
      PC_Next_fetch_5_port, PC_Next_fetch_4_port, PC_Next_fetch_3_port, 
      PC_Next_fetch_2_port, PC_Next_fetch_1_port, PC_Next_fetch_0_port, 
      IRAM_31_port, IRAM_30_port, IRAM_29_port, IRAM_28_port, IRAM_27_port, 
      IRAM_26_port, IRAM_25_port, IRAM_24_port, IRAM_23_port, IRAM_22_port, 
      IRAM_21_port, IRAM_20_port, IRAM_19_port, IRAM_18_port, IRAM_17_port, 
      IRAM_16_port, IRAM_15_port, IRAM_14_port, IRAM_13_port, IRAM_12_port, 
      IRAM_11_port, IRAM_10_port, IRAM_9_port, IRAM_8_port, IRAM_7_port, 
      IRAM_6_port, IRAM_5_port, IRAM_4_port, IRAM_3_port, IRAM_2_port, 
      IRAM_1_port, IRAM_0_port, ADD_RW_4_port, ADD_RW_3_port, ADD_RW_2_port, 
      ADD_RW_1_port, ADD_RW_0_port, RW_R_decode_31_port, RW_R_decode_30_port, 
      RW_R_decode_29_port, RW_R_decode_28_port, RW_R_decode_27_port, 
      RW_R_decode_26_port, RW_R_decode_25_port, RW_R_decode_24_port, 
      RW_R_decode_23_port, RW_R_decode_22_port, RW_R_decode_21_port, 
      RW_R_decode_20_port, RW_R_decode_19_port, RW_R_decode_18_port, 
      RW_R_decode_17_port, RW_R_decode_16_port, RW_R_decode_15_port, 
      RW_R_decode_14_port, RW_R_decode_13_port, RW_R_decode_12_port, 
      RW_R_decode_11_port, RW_R_decode_10_port, RW_R_decode_9_port, 
      RW_R_decode_8_port, RW_R_decode_7_port, RW_R_decode_6_port, 
      RW_R_decode_5_port, RW_R_decode_4_port, RW_R_decode_3_port, 
      RW_R_decode_2_port, RW_R_decode_1_port, RW_R_decode_0_port, 
      RW_I_decode_31_port, RW_I_decode_30_port, RW_I_decode_29_port, 
      RW_I_decode_28_port, RW_I_decode_27_port, RW_I_decode_26_port, 
      RW_I_decode_25_port, RW_I_decode_24_port, RW_I_decode_23_port, 
      RW_I_decode_22_port, RW_I_decode_21_port, RW_I_decode_20_port, 
      RW_I_decode_19_port, RW_I_decode_18_port, RW_I_decode_17_port, 
      RW_I_decode_16_port, RW_I_decode_15_port, RW_I_decode_14_port, 
      RW_I_decode_13_port, RW_I_decode_12_port, RW_I_decode_11_port, 
      RW_I_decode_10_port, RW_I_decode_9_port, RW_I_decode_8_port, 
      RW_I_decode_7_port, RW_I_decode_6_port, RW_I_decode_5_port, 
      RW_I_decode_4_port, RW_I_decode_3_port, RW_I_decode_2_port, 
      RW_I_decode_1_port, RW_I_decode_0_port, J_imm_31_port, J_imm_30_port, 
      J_imm_29_port, J_imm_28_port, J_imm_27_port, J_imm_26_port, J_imm_25_port
      , J_imm_24_port, J_imm_23_port, J_imm_22_port, J_imm_21_port, 
      J_imm_20_port, J_imm_19_port, J_imm_18_port, J_imm_17_port, J_imm_16_port
      , J_imm_15_port, J_imm_14_port, J_imm_13_port, J_imm_12_port, 
      J_imm_11_port, J_imm_10_port, J_imm_9_port, J_imm_8_port, J_imm_7_port, 
      J_imm_6_port, J_imm_5_port, J_imm_4_port, J_imm_3_port, J_imm_2_port, 
      J_imm_1_port, J_imm_0_port, I_imm_31_port, I_imm_30_port, I_imm_29_port, 
      I_imm_28_port, I_imm_27_port, I_imm_26_port, I_imm_25_port, I_imm_24_port
      , I_imm_23_port, I_imm_22_port, I_imm_21_port, I_imm_20_port, 
      I_imm_19_port, I_imm_18_port, I_imm_17_port, I_imm_16_port, I_imm_15_port
      , I_imm_14_port, I_imm_13_port, I_imm_12_port, I_imm_11_port, 
      I_imm_10_port, I_imm_9_port, I_imm_8_port, I_imm_7_port, I_imm_6_port, 
      I_imm_5_port, I_imm_4_port, I_imm_3_port, I_imm_2_port, I_imm_1_port, 
      I_imm_0_port, RD_data_1_31_port, RD_data_1_30_port, RD_data_1_29_port, 
      RD_data_1_28_port, RD_data_1_27_port, RD_data_1_26_port, 
      RD_data_1_25_port, RD_data_1_24_port, RD_data_1_23_port, 
      RD_data_1_22_port, RD_data_1_21_port, RD_data_1_20_port, 
      RD_data_1_19_port, RD_data_1_18_port, RD_data_1_17_port, 
      RD_data_1_16_port, RD_data_1_15_port, RD_data_1_14_port, 
      RD_data_1_13_port, RD_data_1_12_port, RD_data_1_11_port, 
      RD_data_1_10_port, RD_data_1_9_port, RD_data_1_8_port, RD_data_1_7_port, 
      RD_data_1_6_port, RD_data_1_5_port, RD_data_1_4_port, RD_data_1_3_port, 
      RD_data_1_2_port, RD_data_1_1_port, RD_data_1_0_port, RD_data_2_31_port, 
      RD_data_2_30_port, RD_data_2_29_port, RD_data_2_28_port, 
      RD_data_2_27_port, RD_data_2_26_port, RD_data_2_25_port, 
      RD_data_2_24_port, RD_data_2_23_port, RD_data_2_22_port, 
      RD_data_2_21_port, RD_data_2_20_port, RD_data_2_19_port, 
      RD_data_2_18_port, RD_data_2_17_port, RD_data_2_16_port, 
      RD_data_2_15_port, RD_data_2_14_port, RD_data_2_13_port, 
      RD_data_2_12_port, RD_data_2_11_port, RD_data_2_10_port, RD_data_2_9_port
      , RD_data_2_8_port, RD_data_2_7_port, RD_data_2_6_port, RD_data_2_5_port,
      RD_data_2_4_port, RD_data_2_3_port, RD_data_2_2_port, RD_data_2_1_port, 
      RD_data_2_0_port, PC_Next_decode_31_port, PC_Next_decode_30_port, 
      PC_Next_decode_29_port, PC_Next_decode_28_port, PC_Next_decode_27_port, 
      PC_Next_decode_26_port, PC_Next_decode_25_port, PC_Next_decode_24_port, 
      PC_Next_decode_23_port, PC_Next_decode_22_port, PC_Next_decode_21_port, 
      PC_Next_decode_20_port, PC_Next_decode_19_port, PC_Next_decode_18_port, 
      PC_Next_decode_17_port, PC_Next_decode_16_port, PC_Next_decode_15_port, 
      PC_Next_decode_14_port, PC_Next_decode_13_port, PC_Next_decode_12_port, 
      PC_Next_decode_11_port, PC_Next_decode_10_port, PC_Next_decode_9_port, 
      PC_Next_decode_8_port, PC_Next_decode_7_port, PC_Next_decode_6_port, 
      PC_Next_decode_5_port, PC_Next_decode_4_port, PC_Next_decode_3_port, 
      PC_Next_decode_2_port, PC_Next_decode_1_port, PC_Next_decode_0_port, 
      alu_out_31_port, alu_out_30_port, alu_out_29_port, alu_out_28_port, 
      alu_out_27_port, alu_out_26_port, alu_out_25_port, alu_out_24_port, 
      alu_out_23_port, alu_out_22_port, alu_out_21_port, alu_out_20_port, 
      alu_out_19_port, alu_out_18_port, alu_out_17_port, alu_out_16_port, 
      alu_out_15_port, alu_out_14_port, alu_out_13_port, alu_out_12_port, 
      alu_out_11_port, alu_out_10_port, alu_out_9_port, alu_out_8_port, 
      alu_out_7_port, alu_out_6_port, alu_out_5_port, alu_out_4_port, 
      alu_out_3_port, alu_out_2_port, alu_out_1_port, alu_out_0_port, 
      aluR2_to_mem_31_port, aluR2_to_mem_30_port, aluR2_to_mem_29_port, 
      aluR2_to_mem_28_port, aluR2_to_mem_27_port, aluR2_to_mem_26_port, 
      aluR2_to_mem_25_port, aluR2_to_mem_24_port, aluR2_to_mem_23_port, 
      aluR2_to_mem_22_port, aluR2_to_mem_21_port, aluR2_to_mem_20_port, 
      aluR2_to_mem_19_port, aluR2_to_mem_18_port, aluR2_to_mem_17_port, 
      aluR2_to_mem_16_port, aluR2_to_mem_15_port, aluR2_to_mem_14_port, 
      aluR2_to_mem_13_port, aluR2_to_mem_12_port, aluR2_to_mem_11_port, 
      aluR2_to_mem_10_port, aluR2_to_mem_9_port, aluR2_to_mem_8_port, 
      aluR2_to_mem_7_port, aluR2_to_mem_6_port, aluR2_to_mem_5_port, 
      aluR2_to_mem_4_port, aluR2_to_mem_3_port, aluR2_to_mem_2_port, 
      aluR2_to_mem_1_port, aluR2_to_mem_0_port, b_from_ex_to_mem_31_port, 
      b_from_ex_to_mem_30_port, b_from_ex_to_mem_29_port, 
      b_from_ex_to_mem_28_port, b_from_ex_to_mem_27_port, 
      b_from_ex_to_mem_26_port, b_from_ex_to_mem_25_port, 
      b_from_ex_to_mem_24_port, b_from_ex_to_mem_23_port, 
      b_from_ex_to_mem_22_port, b_from_ex_to_mem_21_port, 
      b_from_ex_to_mem_20_port, b_from_ex_to_mem_19_port, 
      b_from_ex_to_mem_18_port, b_from_ex_to_mem_17_port, 
      b_from_ex_to_mem_16_port, b_from_ex_to_mem_15_port, 
      b_from_ex_to_mem_14_port, b_from_ex_to_mem_13_port, 
      b_from_ex_to_mem_12_port, b_from_ex_to_mem_11_port, 
      b_from_ex_to_mem_10_port, b_from_ex_to_mem_9_port, 
      b_from_ex_to_mem_8_port, b_from_ex_to_mem_7_port, b_from_ex_to_mem_6_port
      , b_from_ex_to_mem_5_port, b_from_ex_to_mem_4_port, 
      b_from_ex_to_mem_3_port, b_from_ex_to_mem_2_port, b_from_ex_to_mem_1_port
      , b_from_ex_to_mem_0_port, pc_from_ex_to_mem_31_port, 
      pc_from_ex_to_mem_30_port, pc_from_ex_to_mem_29_port, 
      pc_from_ex_to_mem_28_port, pc_from_ex_to_mem_27_port, 
      pc_from_ex_to_mem_26_port, pc_from_ex_to_mem_25_port, 
      pc_from_ex_to_mem_24_port, pc_from_ex_to_mem_23_port, 
      pc_from_ex_to_mem_22_port, pc_from_ex_to_mem_21_port, 
      pc_from_ex_to_mem_20_port, pc_from_ex_to_mem_19_port, 
      pc_from_ex_to_mem_18_port, pc_from_ex_to_mem_17_port, 
      pc_from_ex_to_mem_16_port, pc_from_ex_to_mem_15_port, 
      pc_from_ex_to_mem_14_port, pc_from_ex_to_mem_13_port, 
      pc_from_ex_to_mem_12_port, pc_from_ex_to_mem_11_port, 
      pc_from_ex_to_mem_10_port, pc_from_ex_to_mem_9_port, 
      pc_from_ex_to_mem_8_port, pc_from_ex_to_mem_7_port, 
      pc_from_ex_to_mem_6_port, pc_from_ex_to_mem_5_port, 
      pc_from_ex_to_mem_4_port, pc_from_ex_to_mem_3_port, 
      pc_from_ex_to_mem_2_port, pc_from_ex_to_mem_1_port, 
      pc_from_ex_to_mem_0_port, rw_from_ex_to_mem_31_port, 
      rw_from_ex_to_mem_30_port, rw_from_ex_to_mem_29_port, 
      rw_from_ex_to_mem_28_port, rw_from_ex_to_mem_27_port, 
      rw_from_ex_to_mem_26_port, rw_from_ex_to_mem_25_port, 
      rw_from_ex_to_mem_24_port, rw_from_ex_to_mem_23_port, 
      rw_from_ex_to_mem_22_port, rw_from_ex_to_mem_21_port, 
      rw_from_ex_to_mem_20_port, rw_from_ex_to_mem_19_port, 
      rw_from_ex_to_mem_18_port, rw_from_ex_to_mem_17_port, 
      rw_from_ex_to_mem_16_port, rw_from_ex_to_mem_15_port, 
      rw_from_ex_to_mem_14_port, rw_from_ex_to_mem_13_port, 
      rw_from_ex_to_mem_12_port, rw_from_ex_to_mem_11_port, 
      rw_from_ex_to_mem_10_port, rw_from_ex_to_mem_9_port, 
      rw_from_ex_to_mem_8_port, rw_from_ex_to_mem_7_port, 
      rw_from_ex_to_mem_6_port, rw_from_ex_to_mem_5_port, 
      rw_from_ex_to_mem_4_port, rw_from_ex_to_mem_3_port, 
      rw_from_ex_to_mem_2_port, rw_from_ex_to_mem_1_port, 
      rw_from_ex_to_mem_0_port, j_from_ex_to_mem_31_port, 
      j_from_ex_to_mem_30_port, j_from_ex_to_mem_29_port, 
      j_from_ex_to_mem_28_port, j_from_ex_to_mem_27_port, 
      j_from_ex_to_mem_26_port, j_from_ex_to_mem_25_port, 
      j_from_ex_to_mem_24_port, j_from_ex_to_mem_23_port, 
      j_from_ex_to_mem_22_port, j_from_ex_to_mem_21_port, 
      j_from_ex_to_mem_20_port, j_from_ex_to_mem_19_port, 
      j_from_ex_to_mem_18_port, j_from_ex_to_mem_17_port, 
      j_from_ex_to_mem_16_port, j_from_ex_to_mem_15_port, 
      j_from_ex_to_mem_14_port, j_from_ex_to_mem_13_port, 
      j_from_ex_to_mem_12_port, j_from_ex_to_mem_11_port, 
      j_from_ex_to_mem_10_port, j_from_ex_to_mem_9_port, 
      j_from_ex_to_mem_8_port, j_from_ex_to_mem_7_port, j_from_ex_to_mem_6_port
      , j_from_ex_to_mem_5_port, j_from_ex_to_mem_4_port, 
      j_from_ex_to_mem_3_port, j_from_ex_to_mem_2_port, j_from_ex_to_mem_1_port
      , j_from_ex_to_mem_0_port, alu_out_mem_31_port, alu_out_mem_30_port, 
      alu_out_mem_29_port, alu_out_mem_28_port, alu_out_mem_27_port, 
      alu_out_mem_26_port, alu_out_mem_25_port, alu_out_mem_24_port, 
      alu_out_mem_23_port, alu_out_mem_22_port, alu_out_mem_21_port, 
      alu_out_mem_20_port, alu_out_mem_19_port, alu_out_mem_18_port, 
      alu_out_mem_17_port, alu_out_mem_16_port, alu_out_mem_15_port, 
      alu_out_mem_14_port, alu_out_mem_13_port, alu_out_mem_12_port, 
      alu_out_mem_11_port, alu_out_mem_10_port, alu_out_mem_9_port, 
      alu_out_mem_8_port, alu_out_mem_7_port, alu_out_mem_6_port, 
      alu_out_mem_5_port, alu_out_mem_4_port, alu_out_mem_3_port, 
      alu_out_mem_2_port, alu_out_mem_1_port, alu_out_mem_0_port, 
      data_from_mem_to_wb_31_port, data_from_mem_to_wb_30_port, 
      data_from_mem_to_wb_29_port, data_from_mem_to_wb_28_port, 
      data_from_mem_to_wb_27_port, data_from_mem_to_wb_26_port, 
      data_from_mem_to_wb_25_port, data_from_mem_to_wb_24_port, 
      data_from_mem_to_wb_23_port, data_from_mem_to_wb_22_port, 
      data_from_mem_to_wb_21_port, data_from_mem_to_wb_20_port, 
      data_from_mem_to_wb_19_port, data_from_mem_to_wb_18_port, 
      data_from_mem_to_wb_17_port, data_from_mem_to_wb_16_port, 
      data_from_mem_to_wb_15_port, data_from_mem_to_wb_14_port, 
      data_from_mem_to_wb_13_port, data_from_mem_to_wb_12_port, 
      data_from_mem_to_wb_11_port, data_from_mem_to_wb_10_port, 
      data_from_mem_to_wb_9_port, data_from_mem_to_wb_8_port, 
      data_from_mem_to_wb_7_port, data_from_mem_to_wb_6_port, 
      data_from_mem_to_wb_5_port, data_from_mem_to_wb_4_port, 
      data_from_mem_to_wb_3_port, data_from_mem_to_wb_2_port, 
      data_from_mem_to_wb_1_port, data_from_mem_to_wb_0_port, n1, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271 : std_logic;

begin
   pipe_out <= ( pipe_out_31_port, pipe_out_30_port, pipe_out_29_port, 
      pipe_out_28_port, pipe_out_27_port, pipe_out_26_port, pipe_out_25_port, 
      pipe_out_24_port, pipe_out_23_port, pipe_out_22_port, pipe_out_21_port, 
      pipe_out_20_port, pipe_out_19_port, pipe_out_18_port, pipe_out_17_port, 
      pipe_out_16_port, pipe_out_15_port, pipe_out_14_port, pipe_out_13_port, 
      pipe_out_12_port, pipe_out_11_port, pipe_out_10_port, pipe_out_9_port, 
      pipe_out_8_port, pipe_out_7_port, pipe_out_6_port, pipe_out_5_port, 
      pipe_out_4_port, pipe_out_3_port, pipe_out_2_port, pipe_out_1_port, 
      pipe_out_0_port );
   
   IFU : fetchUnit_nbit32 port map( Clk => Clk, Rst => n1, en_reg => en_reg_if,
                           PC_branch_jump(31) => pc_from_mem_to_fetch_31_port, 
                           PC_branch_jump(30) => pc_from_mem_to_fetch_30_port, 
                           PC_branch_jump(29) => pc_from_mem_to_fetch_29_port, 
                           PC_branch_jump(28) => pc_from_mem_to_fetch_28_port, 
                           PC_branch_jump(27) => pc_from_mem_to_fetch_27_port, 
                           PC_branch_jump(26) => pc_from_mem_to_fetch_26_port, 
                           PC_branch_jump(25) => pc_from_mem_to_fetch_25_port, 
                           PC_branch_jump(24) => pc_from_mem_to_fetch_24_port, 
                           PC_branch_jump(23) => pc_from_mem_to_fetch_23_port, 
                           PC_branch_jump(22) => pc_from_mem_to_fetch_22_port, 
                           PC_branch_jump(21) => pc_from_mem_to_fetch_21_port, 
                           PC_branch_jump(20) => pc_from_mem_to_fetch_20_port, 
                           PC_branch_jump(19) => pc_from_mem_to_fetch_19_port, 
                           PC_branch_jump(18) => pc_from_mem_to_fetch_18_port, 
                           PC_branch_jump(17) => pc_from_mem_to_fetch_17_port, 
                           PC_branch_jump(16) => pc_from_mem_to_fetch_16_port, 
                           PC_branch_jump(15) => pc_from_mem_to_fetch_15_port, 
                           PC_branch_jump(14) => pc_from_mem_to_fetch_14_port, 
                           PC_branch_jump(13) => pc_from_mem_to_fetch_13_port, 
                           PC_branch_jump(12) => pc_from_mem_to_fetch_12_port, 
                           PC_branch_jump(11) => pc_from_mem_to_fetch_11_port, 
                           PC_branch_jump(10) => pc_from_mem_to_fetch_10_port, 
                           PC_branch_jump(9) => pc_from_mem_to_fetch_9_port, 
                           PC_branch_jump(8) => pc_from_mem_to_fetch_8_port, 
                           PC_branch_jump(7) => pc_from_mem_to_fetch_7_port, 
                           PC_branch_jump(6) => pc_from_mem_to_fetch_6_port, 
                           PC_branch_jump(5) => pc_from_mem_to_fetch_5_port, 
                           PC_branch_jump(4) => pc_from_mem_to_fetch_4_port, 
                           PC_branch_jump(3) => pc_from_mem_to_fetch_3_port, 
                           PC_branch_jump(2) => pc_from_mem_to_fetch_2_port, 
                           PC_branch_jump(1) => pc_from_mem_to_fetch_1_port, 
                           PC_branch_jump(0) => pc_from_mem_to_fetch_0_port, 
                           dout_IRAM(31) => dout_IRAM(31), dout_IRAM(30) => 
                           dout_IRAM(30), dout_IRAM(29) => dout_IRAM(29), 
                           dout_IRAM(28) => dout_IRAM(28), dout_IRAM(27) => 
                           dout_IRAM(27), dout_IRAM(26) => dout_IRAM(26), 
                           dout_IRAM(25) => dout_IRAM(25), dout_IRAM(24) => 
                           dout_IRAM(24), dout_IRAM(23) => dout_IRAM(23), 
                           dout_IRAM(22) => dout_IRAM(22), dout_IRAM(21) => 
                           dout_IRAM(21), dout_IRAM(20) => dout_IRAM(20), 
                           dout_IRAM(19) => dout_IRAM(19), dout_IRAM(18) => 
                           dout_IRAM(18), dout_IRAM(17) => dout_IRAM(17), 
                           dout_IRAM(16) => dout_IRAM(16), dout_IRAM(15) => 
                           dout_IRAM(15), dout_IRAM(14) => dout_IRAM(14), 
                           dout_IRAM(13) => dout_IRAM(13), dout_IRAM(12) => 
                           dout_IRAM(12), dout_IRAM(11) => dout_IRAM(11), 
                           dout_IRAM(10) => dout_IRAM(10), dout_IRAM(9) => 
                           dout_IRAM(9), dout_IRAM(8) => dout_IRAM(8), 
                           dout_IRAM(7) => dout_IRAM(7), dout_IRAM(6) => 
                           dout_IRAM(6), dout_IRAM(5) => dout_IRAM(5), 
                           dout_IRAM(4) => dout_IRAM(4), dout_IRAM(3) => 
                           dout_IRAM(3), dout_IRAM(2) => dout_IRAM(2), 
                           dout_IRAM(1) => dout_IRAM(1), dout_IRAM(0) => 
                           dout_IRAM(0), PC_op => PC_op, PC_Next_out(31) => 
                           PC_Next_fetch_31_port, PC_Next_out(30) => 
                           PC_Next_fetch_30_port, PC_Next_out(29) => 
                           PC_Next_fetch_29_port, PC_Next_out(28) => 
                           PC_Next_fetch_28_port, PC_Next_out(27) => 
                           PC_Next_fetch_27_port, PC_Next_out(26) => 
                           PC_Next_fetch_26_port, PC_Next_out(25) => 
                           PC_Next_fetch_25_port, PC_Next_out(24) => 
                           PC_Next_fetch_24_port, PC_Next_out(23) => 
                           PC_Next_fetch_23_port, PC_Next_out(22) => 
                           PC_Next_fetch_22_port, PC_Next_out(21) => 
                           PC_Next_fetch_21_port, PC_Next_out(20) => 
                           PC_Next_fetch_20_port, PC_Next_out(19) => 
                           PC_Next_fetch_19_port, PC_Next_out(18) => 
                           PC_Next_fetch_18_port, PC_Next_out(17) => 
                           PC_Next_fetch_17_port, PC_Next_out(16) => 
                           PC_Next_fetch_16_port, PC_Next_out(15) => 
                           PC_Next_fetch_15_port, PC_Next_out(14) => 
                           PC_Next_fetch_14_port, PC_Next_out(13) => 
                           PC_Next_fetch_13_port, PC_Next_out(12) => 
                           PC_Next_fetch_12_port, PC_Next_out(11) => 
                           PC_Next_fetch_11_port, PC_Next_out(10) => 
                           PC_Next_fetch_10_port, PC_Next_out(9) => 
                           PC_Next_fetch_9_port, PC_Next_out(8) => 
                           PC_Next_fetch_8_port, PC_Next_out(7) => 
                           PC_Next_fetch_7_port, PC_Next_out(6) => 
                           PC_Next_fetch_6_port, PC_Next_out(5) => 
                           PC_Next_fetch_5_port, PC_Next_out(4) => 
                           PC_Next_fetch_4_port, PC_Next_out(3) => 
                           PC_Next_fetch_3_port, PC_Next_out(2) => 
                           PC_Next_fetch_2_port, PC_Next_out(1) => 
                           PC_Next_fetch_1_port, PC_Next_out(0) => 
                           PC_Next_fetch_0_port, addr_IRAM(31) => addr_IRAM(31)
                           , addr_IRAM(30) => addr_IRAM(30), addr_IRAM(29) => 
                           addr_IRAM(29), addr_IRAM(28) => addr_IRAM(28), 
                           addr_IRAM(27) => addr_IRAM(27), addr_IRAM(26) => 
                           addr_IRAM(26), addr_IRAM(25) => addr_IRAM(25), 
                           addr_IRAM(24) => addr_IRAM(24), addr_IRAM(23) => 
                           addr_IRAM(23), addr_IRAM(22) => addr_IRAM(22), 
                           addr_IRAM(21) => addr_IRAM(21), addr_IRAM(20) => 
                           addr_IRAM(20), addr_IRAM(19) => addr_IRAM(19), 
                           addr_IRAM(18) => addr_IRAM(18), addr_IRAM(17) => 
                           addr_IRAM(17), addr_IRAM(16) => addr_IRAM(16), 
                           addr_IRAM(15) => addr_IRAM(15), addr_IRAM(14) => 
                           addr_IRAM(14), addr_IRAM(13) => addr_IRAM(13), 
                           addr_IRAM(12) => addr_IRAM(12), addr_IRAM(11) => 
                           addr_IRAM(11), addr_IRAM(10) => addr_IRAM(10), 
                           addr_IRAM(9) => addr_IRAM(9), addr_IRAM(8) => 
                           addr_IRAM(8), addr_IRAM(7) => addr_IRAM(7), 
                           addr_IRAM(6) => addr_IRAM(6), addr_IRAM(5) => 
                           addr_IRAM(5), addr_IRAM(4) => addr_IRAM(4), 
                           addr_IRAM(3) => addr_IRAM(3), addr_IRAM(2) => 
                           addr_IRAM(2), addr_IRAM(1) => addr_IRAM(1), 
                           addr_IRAM(0) => addr_IRAM(0), IRAM_reg_out(31) => 
                           IRAM_31_port, IRAM_reg_out(30) => IRAM_30_port, 
                           IRAM_reg_out(29) => IRAM_29_port, IRAM_reg_out(28) 
                           => IRAM_28_port, IRAM_reg_out(27) => IRAM_27_port, 
                           IRAM_reg_out(26) => IRAM_26_port, IRAM_reg_out(25) 
                           => IRAM_25_port, IRAM_reg_out(24) => IRAM_24_port, 
                           IRAM_reg_out(23) => IRAM_23_port, IRAM_reg_out(22) 
                           => IRAM_22_port, IRAM_reg_out(21) => IRAM_21_port, 
                           IRAM_reg_out(20) => IRAM_20_port, IRAM_reg_out(19) 
                           => IRAM_19_port, IRAM_reg_out(18) => IRAM_18_port, 
                           IRAM_reg_out(17) => IRAM_17_port, IRAM_reg_out(16) 
                           => IRAM_16_port, IRAM_reg_out(15) => IRAM_15_port, 
                           IRAM_reg_out(14) => IRAM_14_port, IRAM_reg_out(13) 
                           => IRAM_13_port, IRAM_reg_out(12) => IRAM_12_port, 
                           IRAM_reg_out(11) => IRAM_11_port, IRAM_reg_out(10) 
                           => IRAM_10_port, IRAM_reg_out(9) => IRAM_9_port, 
                           IRAM_reg_out(8) => IRAM_8_port, IRAM_reg_out(7) => 
                           IRAM_7_port, IRAM_reg_out(6) => IRAM_6_port, 
                           IRAM_reg_out(5) => IRAM_5_port, IRAM_reg_out(4) => 
                           IRAM_4_port, IRAM_reg_out(3) => IRAM_3_port, 
                           IRAM_reg_out(2) => IRAM_2_port, IRAM_reg_out(1) => 
                           IRAM_1_port, IRAM_reg_out(0) => IRAM_0_port);
   IDU : decodeUnit_nbit32 port map( Clk => Clk, Rst => n1, en_reg => en_reg_id
                           , RD1 => RD1, RD2 => RD2, IRAM_instr(31) => 
                           IRAM_31_port, IRAM_instr(30) => IRAM_30_port, 
                           IRAM_instr(29) => IRAM_29_port, IRAM_instr(28) => 
                           IRAM_28_port, IRAM_instr(27) => IRAM_27_port, 
                           IRAM_instr(26) => IRAM_26_port, IRAM_instr(25) => 
                           IRAM_25_port, IRAM_instr(24) => IRAM_24_port, 
                           IRAM_instr(23) => IRAM_23_port, IRAM_instr(22) => 
                           IRAM_22_port, IRAM_instr(21) => IRAM_21_port, 
                           IRAM_instr(20) => IRAM_20_port, IRAM_instr(19) => 
                           IRAM_19_port, IRAM_instr(18) => IRAM_18_port, 
                           IRAM_instr(17) => IRAM_17_port, IRAM_instr(16) => 
                           IRAM_16_port, IRAM_instr(15) => IRAM_15_port, 
                           IRAM_instr(14) => IRAM_14_port, IRAM_instr(13) => 
                           IRAM_13_port, IRAM_instr(12) => IRAM_12_port, 
                           IRAM_instr(11) => IRAM_11_port, IRAM_instr(10) => 
                           IRAM_10_port, IRAM_instr(9) => IRAM_9_port, 
                           IRAM_instr(8) => IRAM_8_port, IRAM_instr(7) => 
                           IRAM_7_port, IRAM_instr(6) => IRAM_6_port, 
                           IRAM_instr(5) => IRAM_5_port, IRAM_instr(4) => 
                           IRAM_4_port, IRAM_instr(3) => IRAM_3_port, 
                           IRAM_instr(2) => IRAM_2_port, IRAM_instr(1) => 
                           IRAM_1_port, IRAM_instr(0) => IRAM_0_port, 
                           PC_Next(31) => PC_Next_fetch_31_port, PC_Next(30) =>
                           PC_Next_fetch_30_port, PC_Next(29) => 
                           PC_Next_fetch_29_port, PC_Next(28) => 
                           PC_Next_fetch_28_port, PC_Next(27) => 
                           PC_Next_fetch_27_port, PC_Next(26) => 
                           PC_Next_fetch_26_port, PC_Next(25) => 
                           PC_Next_fetch_25_port, PC_Next(24) => 
                           PC_Next_fetch_24_port, PC_Next(23) => 
                           PC_Next_fetch_23_port, PC_Next(22) => 
                           PC_Next_fetch_22_port, PC_Next(21) => 
                           PC_Next_fetch_21_port, PC_Next(20) => 
                           PC_Next_fetch_20_port, PC_Next(19) => 
                           PC_Next_fetch_19_port, PC_Next(18) => 
                           PC_Next_fetch_18_port, PC_Next(17) => 
                           PC_Next_fetch_17_port, PC_Next(16) => 
                           PC_Next_fetch_16_port, PC_Next(15) => 
                           PC_Next_fetch_15_port, PC_Next(14) => 
                           PC_Next_fetch_14_port, PC_Next(13) => 
                           PC_Next_fetch_13_port, PC_Next(12) => 
                           PC_Next_fetch_12_port, PC_Next(11) => 
                           PC_Next_fetch_11_port, PC_Next(10) => 
                           PC_Next_fetch_10_port, PC_Next(9) => 
                           PC_Next_fetch_9_port, PC_Next(8) => 
                           PC_Next_fetch_8_port, PC_Next(7) => 
                           PC_Next_fetch_7_port, PC_Next(6) => 
                           PC_Next_fetch_6_port, PC_Next(5) => 
                           PC_Next_fetch_5_port, PC_Next(4) => 
                           PC_Next_fetch_4_port, PC_Next(3) => 
                           PC_Next_fetch_3_port, PC_Next(2) => 
                           PC_Next_fetch_2_port, PC_Next(1) => 
                           PC_Next_fetch_1_port, PC_Next(0) => 
                           PC_Next_fetch_0_port, WR => WR, ADD_RW(4) => 
                           ADD_RW_4_port, ADD_RW(3) => ADD_RW_3_port, ADD_RW(2)
                           => ADD_RW_2_port, ADD_RW(1) => ADD_RW_1_port, 
                           ADD_RW(0) => ADD_RW_0_port, DATA_RW(31) => 
                           pipe_out_31_port, DATA_RW(30) => pipe_out_30_port, 
                           DATA_RW(29) => pipe_out_29_port, DATA_RW(28) => 
                           pipe_out_28_port, DATA_RW(27) => pipe_out_27_port, 
                           DATA_RW(26) => pipe_out_26_port, DATA_RW(25) => 
                           pipe_out_25_port, DATA_RW(24) => pipe_out_24_port, 
                           DATA_RW(23) => pipe_out_23_port, DATA_RW(22) => 
                           pipe_out_22_port, DATA_RW(21) => pipe_out_21_port, 
                           DATA_RW(20) => pipe_out_20_port, DATA_RW(19) => 
                           pipe_out_19_port, DATA_RW(18) => pipe_out_18_port, 
                           DATA_RW(17) => pipe_out_17_port, DATA_RW(16) => 
                           pipe_out_16_port, DATA_RW(15) => pipe_out_15_port, 
                           DATA_RW(14) => pipe_out_14_port, DATA_RW(13) => 
                           pipe_out_13_port, DATA_RW(12) => pipe_out_12_port, 
                           DATA_RW(11) => pipe_out_11_port, DATA_RW(10) => 
                           pipe_out_10_port, DATA_RW(9) => pipe_out_9_port, 
                           DATA_RW(8) => pipe_out_8_port, DATA_RW(7) => 
                           pipe_out_7_port, DATA_RW(6) => pipe_out_6_port, 
                           DATA_RW(5) => pipe_out_5_port, DATA_RW(4) => 
                           pipe_out_4_port, DATA_RW(3) => pipe_out_3_port, 
                           DATA_RW(2) => pipe_out_2_port, DATA_RW(1) => 
                           pipe_out_1_port, DATA_RW(0) => pipe_out_0_port, 
                           RW_R_out(31) => RW_R_decode_31_port, RW_R_out(30) =>
                           RW_R_decode_30_port, RW_R_out(29) => 
                           RW_R_decode_29_port, RW_R_out(28) => 
                           RW_R_decode_28_port, RW_R_out(27) => 
                           RW_R_decode_27_port, RW_R_out(26) => 
                           RW_R_decode_26_port, RW_R_out(25) => 
                           RW_R_decode_25_port, RW_R_out(24) => 
                           RW_R_decode_24_port, RW_R_out(23) => 
                           RW_R_decode_23_port, RW_R_out(22) => 
                           RW_R_decode_22_port, RW_R_out(21) => 
                           RW_R_decode_21_port, RW_R_out(20) => 
                           RW_R_decode_20_port, RW_R_out(19) => 
                           RW_R_decode_19_port, RW_R_out(18) => 
                           RW_R_decode_18_port, RW_R_out(17) => 
                           RW_R_decode_17_port, RW_R_out(16) => 
                           RW_R_decode_16_port, RW_R_out(15) => 
                           RW_R_decode_15_port, RW_R_out(14) => 
                           RW_R_decode_14_port, RW_R_out(13) => 
                           RW_R_decode_13_port, RW_R_out(12) => 
                           RW_R_decode_12_port, RW_R_out(11) => 
                           RW_R_decode_11_port, RW_R_out(10) => 
                           RW_R_decode_10_port, RW_R_out(9) => 
                           RW_R_decode_9_port, RW_R_out(8) => 
                           RW_R_decode_8_port, RW_R_out(7) => 
                           RW_R_decode_7_port, RW_R_out(6) => 
                           RW_R_decode_6_port, RW_R_out(5) => 
                           RW_R_decode_5_port, RW_R_out(4) => 
                           RW_R_decode_4_port, RW_R_out(3) => 
                           RW_R_decode_3_port, RW_R_out(2) => 
                           RW_R_decode_2_port, RW_R_out(1) => 
                           RW_R_decode_1_port, RW_R_out(0) => 
                           RW_R_decode_0_port, RW_I_out(31) => 
                           RW_I_decode_31_port, RW_I_out(30) => 
                           RW_I_decode_30_port, RW_I_out(29) => 
                           RW_I_decode_29_port, RW_I_out(28) => 
                           RW_I_decode_28_port, RW_I_out(27) => 
                           RW_I_decode_27_port, RW_I_out(26) => 
                           RW_I_decode_26_port, RW_I_out(25) => 
                           RW_I_decode_25_port, RW_I_out(24) => 
                           RW_I_decode_24_port, RW_I_out(23) => 
                           RW_I_decode_23_port, RW_I_out(22) => 
                           RW_I_decode_22_port, RW_I_out(21) => 
                           RW_I_decode_21_port, RW_I_out(20) => 
                           RW_I_decode_20_port, RW_I_out(19) => 
                           RW_I_decode_19_port, RW_I_out(18) => 
                           RW_I_decode_18_port, RW_I_out(17) => 
                           RW_I_decode_17_port, RW_I_out(16) => 
                           RW_I_decode_16_port, RW_I_out(15) => 
                           RW_I_decode_15_port, RW_I_out(14) => 
                           RW_I_decode_14_port, RW_I_out(13) => 
                           RW_I_decode_13_port, RW_I_out(12) => 
                           RW_I_decode_12_port, RW_I_out(11) => 
                           RW_I_decode_11_port, RW_I_out(10) => 
                           RW_I_decode_10_port, RW_I_out(9) => 
                           RW_I_decode_9_port, RW_I_out(8) => 
                           RW_I_decode_8_port, RW_I_out(7) => 
                           RW_I_decode_7_port, RW_I_out(6) => 
                           RW_I_decode_6_port, RW_I_out(5) => 
                           RW_I_decode_5_port, RW_I_out(4) => 
                           RW_I_decode_4_port, RW_I_out(3) => 
                           RW_I_decode_3_port, RW_I_out(2) => 
                           RW_I_decode_2_port, RW_I_out(1) => 
                           RW_I_decode_1_port, RW_I_out(0) => 
                           RW_I_decode_0_port, Jump_address(31) => 
                           J_imm_31_port, Jump_address(30) => J_imm_30_port, 
                           Jump_address(29) => J_imm_29_port, Jump_address(28) 
                           => J_imm_28_port, Jump_address(27) => J_imm_27_port,
                           Jump_address(26) => J_imm_26_port, Jump_address(25) 
                           => J_imm_25_port, Jump_address(24) => J_imm_24_port,
                           Jump_address(23) => J_imm_23_port, Jump_address(22) 
                           => J_imm_22_port, Jump_address(21) => J_imm_21_port,
                           Jump_address(20) => J_imm_20_port, Jump_address(19) 
                           => J_imm_19_port, Jump_address(18) => J_imm_18_port,
                           Jump_address(17) => J_imm_17_port, Jump_address(16) 
                           => J_imm_16_port, Jump_address(15) => J_imm_15_port,
                           Jump_address(14) => J_imm_14_port, Jump_address(13) 
                           => J_imm_13_port, Jump_address(12) => J_imm_12_port,
                           Jump_address(11) => J_imm_11_port, Jump_address(10) 
                           => J_imm_10_port, Jump_address(9) => J_imm_9_port, 
                           Jump_address(8) => J_imm_8_port, Jump_address(7) => 
                           J_imm_7_port, Jump_address(6) => J_imm_6_port, 
                           Jump_address(5) => J_imm_5_port, Jump_address(4) => 
                           J_imm_4_port, Jump_address(3) => J_imm_3_port, 
                           Jump_address(2) => J_imm_2_port, Jump_address(1) => 
                           J_imm_1_port, Jump_address(0) => J_imm_0_port, 
                           I_immediate_ext_out(31) => I_imm_31_port, 
                           I_immediate_ext_out(30) => I_imm_30_port, 
                           I_immediate_ext_out(29) => I_imm_29_port, 
                           I_immediate_ext_out(28) => I_imm_28_port, 
                           I_immediate_ext_out(27) => I_imm_27_port, 
                           I_immediate_ext_out(26) => I_imm_26_port, 
                           I_immediate_ext_out(25) => I_imm_25_port, 
                           I_immediate_ext_out(24) => I_imm_24_port, 
                           I_immediate_ext_out(23) => I_imm_23_port, 
                           I_immediate_ext_out(22) => I_imm_22_port, 
                           I_immediate_ext_out(21) => I_imm_21_port, 
                           I_immediate_ext_out(20) => I_imm_20_port, 
                           I_immediate_ext_out(19) => I_imm_19_port, 
                           I_immediate_ext_out(18) => I_imm_18_port, 
                           I_immediate_ext_out(17) => I_imm_17_port, 
                           I_immediate_ext_out(16) => I_imm_16_port, 
                           I_immediate_ext_out(15) => I_imm_15_port, 
                           I_immediate_ext_out(14) => I_imm_14_port, 
                           I_immediate_ext_out(13) => I_imm_13_port, 
                           I_immediate_ext_out(12) => I_imm_12_port, 
                           I_immediate_ext_out(11) => I_imm_11_port, 
                           I_immediate_ext_out(10) => I_imm_10_port, 
                           I_immediate_ext_out(9) => I_imm_9_port, 
                           I_immediate_ext_out(8) => I_imm_8_port, 
                           I_immediate_ext_out(7) => I_imm_7_port, 
                           I_immediate_ext_out(6) => I_imm_6_port, 
                           I_immediate_ext_out(5) => I_imm_5_port, 
                           I_immediate_ext_out(4) => I_imm_4_port, 
                           I_immediate_ext_out(3) => I_imm_3_port, 
                           I_immediate_ext_out(2) => I_imm_2_port, 
                           I_immediate_ext_out(1) => I_imm_1_port, 
                           I_immediate_ext_out(0) => I_imm_0_port, 
                           RD_data_1_out(31) => RD_data_1_31_port, 
                           RD_data_1_out(30) => RD_data_1_30_port, 
                           RD_data_1_out(29) => RD_data_1_29_port, 
                           RD_data_1_out(28) => RD_data_1_28_port, 
                           RD_data_1_out(27) => RD_data_1_27_port, 
                           RD_data_1_out(26) => RD_data_1_26_port, 
                           RD_data_1_out(25) => RD_data_1_25_port, 
                           RD_data_1_out(24) => RD_data_1_24_port, 
                           RD_data_1_out(23) => RD_data_1_23_port, 
                           RD_data_1_out(22) => RD_data_1_22_port, 
                           RD_data_1_out(21) => RD_data_1_21_port, 
                           RD_data_1_out(20) => RD_data_1_20_port, 
                           RD_data_1_out(19) => RD_data_1_19_port, 
                           RD_data_1_out(18) => RD_data_1_18_port, 
                           RD_data_1_out(17) => RD_data_1_17_port, 
                           RD_data_1_out(16) => RD_data_1_16_port, 
                           RD_data_1_out(15) => RD_data_1_15_port, 
                           RD_data_1_out(14) => RD_data_1_14_port, 
                           RD_data_1_out(13) => RD_data_1_13_port, 
                           RD_data_1_out(12) => RD_data_1_12_port, 
                           RD_data_1_out(11) => RD_data_1_11_port, 
                           RD_data_1_out(10) => RD_data_1_10_port, 
                           RD_data_1_out(9) => RD_data_1_9_port, 
                           RD_data_1_out(8) => RD_data_1_8_port, 
                           RD_data_1_out(7) => RD_data_1_7_port, 
                           RD_data_1_out(6) => RD_data_1_6_port, 
                           RD_data_1_out(5) => RD_data_1_5_port, 
                           RD_data_1_out(4) => RD_data_1_4_port, 
                           RD_data_1_out(3) => RD_data_1_3_port, 
                           RD_data_1_out(2) => RD_data_1_2_port, 
                           RD_data_1_out(1) => RD_data_1_1_port, 
                           RD_data_1_out(0) => RD_data_1_0_port, 
                           RD_data_2_out(31) => RD_data_2_31_port, 
                           RD_data_2_out(30) => RD_data_2_30_port, 
                           RD_data_2_out(29) => RD_data_2_29_port, 
                           RD_data_2_out(28) => RD_data_2_28_port, 
                           RD_data_2_out(27) => RD_data_2_27_port, 
                           RD_data_2_out(26) => RD_data_2_26_port, 
                           RD_data_2_out(25) => RD_data_2_25_port, 
                           RD_data_2_out(24) => RD_data_2_24_port, 
                           RD_data_2_out(23) => RD_data_2_23_port, 
                           RD_data_2_out(22) => RD_data_2_22_port, 
                           RD_data_2_out(21) => RD_data_2_21_port, 
                           RD_data_2_out(20) => RD_data_2_20_port, 
                           RD_data_2_out(19) => RD_data_2_19_port, 
                           RD_data_2_out(18) => RD_data_2_18_port, 
                           RD_data_2_out(17) => RD_data_2_17_port, 
                           RD_data_2_out(16) => RD_data_2_16_port, 
                           RD_data_2_out(15) => RD_data_2_15_port, 
                           RD_data_2_out(14) => RD_data_2_14_port, 
                           RD_data_2_out(13) => RD_data_2_13_port, 
                           RD_data_2_out(12) => RD_data_2_12_port, 
                           RD_data_2_out(11) => RD_data_2_11_port, 
                           RD_data_2_out(10) => RD_data_2_10_port, 
                           RD_data_2_out(9) => RD_data_2_9_port, 
                           RD_data_2_out(8) => RD_data_2_8_port, 
                           RD_data_2_out(7) => RD_data_2_7_port, 
                           RD_data_2_out(6) => RD_data_2_6_port, 
                           RD_data_2_out(5) => RD_data_2_5_port, 
                           RD_data_2_out(4) => RD_data_2_4_port, 
                           RD_data_2_out(3) => RD_data_2_3_port, 
                           RD_data_2_out(2) => RD_data_2_2_port, 
                           RD_data_2_out(1) => RD_data_2_1_port, 
                           RD_data_2_out(0) => RD_data_2_0_port, 
                           PC_Next_out(31) => PC_Next_decode_31_port, 
                           PC_Next_out(30) => PC_Next_decode_30_port, 
                           PC_Next_out(29) => PC_Next_decode_29_port, 
                           PC_Next_out(28) => PC_Next_decode_28_port, 
                           PC_Next_out(27) => PC_Next_decode_27_port, 
                           PC_Next_out(26) => PC_Next_decode_26_port, 
                           PC_Next_out(25) => PC_Next_decode_25_port, 
                           PC_Next_out(24) => PC_Next_decode_24_port, 
                           PC_Next_out(23) => PC_Next_decode_23_port, 
                           PC_Next_out(22) => PC_Next_decode_22_port, 
                           PC_Next_out(21) => PC_Next_decode_21_port, 
                           PC_Next_out(20) => PC_Next_decode_20_port, 
                           PC_Next_out(19) => PC_Next_decode_19_port, 
                           PC_Next_out(18) => PC_Next_decode_18_port, 
                           PC_Next_out(17) => PC_Next_decode_17_port, 
                           PC_Next_out(16) => PC_Next_decode_16_port, 
                           PC_Next_out(15) => PC_Next_decode_15_port, 
                           PC_Next_out(14) => PC_Next_decode_14_port, 
                           PC_Next_out(13) => PC_Next_decode_13_port, 
                           PC_Next_out(12) => PC_Next_decode_12_port, 
                           PC_Next_out(11) => PC_Next_decode_11_port, 
                           PC_Next_out(10) => PC_Next_decode_10_port, 
                           PC_Next_out(9) => PC_Next_decode_9_port, 
                           PC_Next_out(8) => PC_Next_decode_8_port, 
                           PC_Next_out(7) => PC_Next_decode_7_port, 
                           PC_Next_out(6) => PC_Next_decode_6_port, 
                           PC_Next_out(5) => PC_Next_decode_5_port, 
                           PC_Next_out(4) => PC_Next_decode_4_port, 
                           PC_Next_out(3) => PC_Next_decode_3_port, 
                           PC_Next_out(2) => PC_Next_decode_2_port, 
                           PC_Next_out(1) => PC_Next_decode_1_port, 
                           PC_Next_out(0) => PC_Next_decode_0_port, Opcode(5) 
                           => Opcode(5), Opcode(4) => Opcode(4), Opcode(3) => 
                           Opcode(3), Opcode(2) => Opcode(2), Opcode(1) => 
                           Opcode(1), Opcode(0) => Opcode(0), Func(10) => 
                           Func(10), Func(9) => Func(9), Func(8) => Func(8), 
                           Func(7) => Func(7), Func(6) => Func(6), Func(5) => 
                           Func(5), Func(4) => Func(4), Func(3) => Func(3), 
                           Func(2) => Func(2), Func(1) => Func(1), Func(0) => 
                           Func(0));
   EXE : executionUnit_nbit32 port map( r1(31) => RD_data_1_31_port, r1(30) => 
                           RD_data_1_30_port, r1(29) => RD_data_1_29_port, 
                           r1(28) => RD_data_1_28_port, r1(27) => 
                           RD_data_1_27_port, r1(26) => RD_data_1_26_port, 
                           r1(25) => RD_data_1_25_port, r1(24) => 
                           RD_data_1_24_port, r1(23) => RD_data_1_23_port, 
                           r1(22) => RD_data_1_22_port, r1(21) => 
                           RD_data_1_21_port, r1(20) => RD_data_1_20_port, 
                           r1(19) => RD_data_1_19_port, r1(18) => 
                           RD_data_1_18_port, r1(17) => RD_data_1_17_port, 
                           r1(16) => RD_data_1_16_port, r1(15) => 
                           RD_data_1_15_port, r1(14) => RD_data_1_14_port, 
                           r1(13) => RD_data_1_13_port, r1(12) => 
                           RD_data_1_12_port, r1(11) => RD_data_1_11_port, 
                           r1(10) => RD_data_1_10_port, r1(9) => 
                           RD_data_1_9_port, r1(8) => RD_data_1_8_port, r1(7) 
                           => RD_data_1_7_port, r1(6) => RD_data_1_6_port, 
                           r1(5) => RD_data_1_5_port, r1(4) => RD_data_1_4_port
                           , r1(3) => RD_data_1_3_port, r1(2) => 
                           RD_data_1_2_port, r1(1) => RD_data_1_1_port, r1(0) 
                           => RD_data_1_0_port, r2(31) => RD_data_2_31_port, 
                           r2(30) => RD_data_2_30_port, r2(29) => 
                           RD_data_2_29_port, r2(28) => RD_data_2_28_port, 
                           r2(27) => RD_data_2_27_port, r2(26) => 
                           RD_data_2_26_port, r2(25) => RD_data_2_25_port, 
                           r2(24) => RD_data_2_24_port, r2(23) => 
                           RD_data_2_23_port, r2(22) => RD_data_2_22_port, 
                           r2(21) => RD_data_2_21_port, r2(20) => 
                           RD_data_2_20_port, r2(19) => RD_data_2_19_port, 
                           r2(18) => RD_data_2_18_port, r2(17) => 
                           RD_data_2_17_port, r2(16) => RD_data_2_16_port, 
                           r2(15) => RD_data_2_15_port, r2(14) => 
                           RD_data_2_14_port, r2(13) => RD_data_2_13_port, 
                           r2(12) => RD_data_2_12_port, r2(11) => 
                           RD_data_2_11_port, r2(10) => RD_data_2_10_port, 
                           r2(9) => RD_data_2_9_port, r2(8) => RD_data_2_8_port
                           , r2(7) => RD_data_2_7_port, r2(6) => 
                           RD_data_2_6_port, r2(5) => RD_data_2_5_port, r2(4) 
                           => RD_data_2_4_port, r2(3) => RD_data_2_3_port, 
                           r2(2) => RD_data_2_2_port, r2(1) => RD_data_2_1_port
                           , r2(0) => RD_data_2_0_port, imm(31) => 
                           I_imm_31_port, imm(30) => I_imm_30_port, imm(29) => 
                           I_imm_29_port, imm(28) => I_imm_28_port, imm(27) => 
                           I_imm_27_port, imm(26) => I_imm_26_port, imm(25) => 
                           I_imm_25_port, imm(24) => I_imm_24_port, imm(23) => 
                           I_imm_23_port, imm(22) => I_imm_22_port, imm(21) => 
                           I_imm_21_port, imm(20) => I_imm_20_port, imm(19) => 
                           I_imm_19_port, imm(18) => I_imm_18_port, imm(17) => 
                           I_imm_17_port, imm(16) => I_imm_16_port, imm(15) => 
                           I_imm_15_port, imm(14) => I_imm_14_port, imm(13) => 
                           I_imm_13_port, imm(12) => I_imm_12_port, imm(11) => 
                           I_imm_11_port, imm(10) => I_imm_10_port, imm(9) => 
                           I_imm_9_port, imm(8) => I_imm_8_port, imm(7) => 
                           I_imm_7_port, imm(6) => I_imm_6_port, imm(5) => 
                           I_imm_5_port, imm(4) => I_imm_4_port, imm(3) => 
                           I_imm_3_port, imm(2) => I_imm_2_port, imm(1) => 
                           I_imm_1_port, imm(0) => I_imm_0_port, j_lab(31) => 
                           J_imm_31_port, j_lab(30) => J_imm_30_port, j_lab(29)
                           => J_imm_29_port, j_lab(28) => J_imm_28_port, 
                           j_lab(27) => J_imm_27_port, j_lab(26) => 
                           J_imm_26_port, j_lab(25) => J_imm_25_port, j_lab(24)
                           => J_imm_24_port, j_lab(23) => J_imm_23_port, 
                           j_lab(22) => J_imm_22_port, j_lab(21) => 
                           J_imm_21_port, j_lab(20) => J_imm_20_port, j_lab(19)
                           => J_imm_19_port, j_lab(18) => J_imm_18_port, 
                           j_lab(17) => J_imm_17_port, j_lab(16) => 
                           J_imm_16_port, j_lab(15) => J_imm_15_port, j_lab(14)
                           => J_imm_14_port, j_lab(13) => J_imm_13_port, 
                           j_lab(12) => J_imm_12_port, j_lab(11) => 
                           J_imm_11_port, j_lab(10) => J_imm_10_port, j_lab(9) 
                           => J_imm_9_port, j_lab(8) => J_imm_8_port, j_lab(7) 
                           => J_imm_7_port, j_lab(6) => J_imm_6_port, j_lab(5) 
                           => J_imm_5_port, j_lab(4) => J_imm_4_port, j_lab(3) 
                           => J_imm_3_port, j_lab(2) => J_imm_2_port, j_lab(1) 
                           => J_imm_1_port, j_lab(0) => J_imm_0_port, pc(31) =>
                           PC_Next_decode_31_port, pc(30) => 
                           PC_Next_decode_30_port, pc(29) => 
                           PC_Next_decode_29_port, pc(28) => 
                           PC_Next_decode_28_port, pc(27) => 
                           PC_Next_decode_27_port, pc(26) => 
                           PC_Next_decode_26_port, pc(25) => 
                           PC_Next_decode_25_port, pc(24) => 
                           PC_Next_decode_24_port, pc(23) => 
                           PC_Next_decode_23_port, pc(22) => 
                           PC_Next_decode_22_port, pc(21) => 
                           PC_Next_decode_21_port, pc(20) => 
                           PC_Next_decode_20_port, pc(19) => 
                           PC_Next_decode_19_port, pc(18) => 
                           PC_Next_decode_18_port, pc(17) => 
                           PC_Next_decode_17_port, pc(16) => 
                           PC_Next_decode_16_port, pc(15) => 
                           PC_Next_decode_15_port, pc(14) => 
                           PC_Next_decode_14_port, pc(13) => 
                           PC_Next_decode_13_port, pc(12) => 
                           PC_Next_decode_12_port, pc(11) => 
                           PC_Next_decode_11_port, pc(10) => 
                           PC_Next_decode_10_port, pc(9) => 
                           PC_Next_decode_9_port, pc(8) => 
                           PC_Next_decode_8_port, pc(7) => 
                           PC_Next_decode_7_port, pc(6) => 
                           PC_Next_decode_6_port, pc(5) => 
                           PC_Next_decode_5_port, pc(4) => 
                           PC_Next_decode_4_port, pc(3) => 
                           PC_Next_decode_3_port, pc(2) => 
                           PC_Next_decode_2_port, pc(1) => 
                           PC_Next_decode_1_port, pc(0) => 
                           PC_Next_decode_0_port, RW_R(31) => 
                           RW_R_decode_31_port, RW_R(30) => RW_R_decode_30_port
                           , RW_R(29) => RW_R_decode_29_port, RW_R(28) => 
                           RW_R_decode_28_port, RW_R(27) => RW_R_decode_27_port
                           , RW_R(26) => RW_R_decode_26_port, RW_R(25) => 
                           RW_R_decode_25_port, RW_R(24) => RW_R_decode_24_port
                           , RW_R(23) => RW_R_decode_23_port, RW_R(22) => 
                           RW_R_decode_22_port, RW_R(21) => RW_R_decode_21_port
                           , RW_R(20) => RW_R_decode_20_port, RW_R(19) => 
                           RW_R_decode_19_port, RW_R(18) => RW_R_decode_18_port
                           , RW_R(17) => RW_R_decode_17_port, RW_R(16) => 
                           RW_R_decode_16_port, RW_R(15) => RW_R_decode_15_port
                           , RW_R(14) => RW_R_decode_14_port, RW_R(13) => 
                           RW_R_decode_13_port, RW_R(12) => RW_R_decode_12_port
                           , RW_R(11) => RW_R_decode_11_port, RW_R(10) => 
                           RW_R_decode_10_port, RW_R(9) => RW_R_decode_9_port, 
                           RW_R(8) => RW_R_decode_8_port, RW_R(7) => 
                           RW_R_decode_7_port, RW_R(6) => RW_R_decode_6_port, 
                           RW_R(5) => RW_R_decode_5_port, RW_R(4) => 
                           RW_R_decode_4_port, RW_R(3) => RW_R_decode_3_port, 
                           RW_R(2) => RW_R_decode_2_port, RW_R(1) => 
                           RW_R_decode_1_port, RW_R(0) => RW_R_decode_0_port, 
                           RW_I(31) => RW_I_decode_31_port, RW_I(30) => 
                           RW_I_decode_30_port, RW_I(29) => RW_I_decode_29_port
                           , RW_I(28) => RW_I_decode_28_port, RW_I(27) => 
                           RW_I_decode_27_port, RW_I(26) => RW_I_decode_26_port
                           , RW_I(25) => RW_I_decode_25_port, RW_I(24) => 
                           RW_I_decode_24_port, RW_I(23) => RW_I_decode_23_port
                           , RW_I(22) => RW_I_decode_22_port, RW_I(21) => 
                           RW_I_decode_21_port, RW_I(20) => RW_I_decode_20_port
                           , RW_I(19) => RW_I_decode_19_port, RW_I(18) => 
                           RW_I_decode_18_port, RW_I(17) => RW_I_decode_17_port
                           , RW_I(16) => RW_I_decode_16_port, RW_I(15) => 
                           RW_I_decode_15_port, RW_I(14) => RW_I_decode_14_port
                           , RW_I(13) => RW_I_decode_13_port, RW_I(12) => 
                           RW_I_decode_12_port, RW_I(11) => RW_I_decode_11_port
                           , RW_I(10) => RW_I_decode_10_port, RW_I(9) => 
                           RW_I_decode_9_port, RW_I(8) => RW_I_decode_8_port, 
                           RW_I(7) => RW_I_decode_7_port, RW_I(6) => 
                           RW_I_decode_6_port, RW_I(5) => RW_I_decode_5_port, 
                           RW_I(4) => RW_I_decode_4_port, RW_I(3) => 
                           RW_I_decode_3_port, RW_I(2) => RW_I_decode_2_port, 
                           RW_I(1) => RW_I_decode_1_port, RW_I(0) => 
                           RW_I_decode_0_port, s2 => sel_ex, s3 => sel_mux_rw, 
                           rst => n1, clk => Clk, en_reg => en_reg_ex, 
                           alu_sel(3) => alu_sel(3), alu_sel(2) => alu_sel(2), 
                           alu_sel(1) => alu_sel(1), alu_sel(0) => alu_sel(0), 
                           alu_out(31) => alu_out_31_port, alu_out(30) => 
                           alu_out_30_port, alu_out(29) => alu_out_29_port, 
                           alu_out(28) => alu_out_28_port, alu_out(27) => 
                           alu_out_27_port, alu_out(26) => alu_out_26_port, 
                           alu_out(25) => alu_out_25_port, alu_out(24) => 
                           alu_out_24_port, alu_out(23) => alu_out_23_port, 
                           alu_out(22) => alu_out_22_port, alu_out(21) => 
                           alu_out_21_port, alu_out(20) => alu_out_20_port, 
                           alu_out(19) => alu_out_19_port, alu_out(18) => 
                           alu_out_18_port, alu_out(17) => alu_out_17_port, 
                           alu_out(16) => alu_out_16_port, alu_out(15) => 
                           alu_out_15_port, alu_out(14) => alu_out_14_port, 
                           alu_out(13) => alu_out_13_port, alu_out(12) => 
                           alu_out_12_port, alu_out(11) => alu_out_11_port, 
                           alu_out(10) => alu_out_10_port, alu_out(9) => 
                           alu_out_9_port, alu_out(8) => alu_out_8_port, 
                           alu_out(7) => alu_out_7_port, alu_out(6) => 
                           alu_out_6_port, alu_out(5) => alu_out_5_port, 
                           alu_out(4) => alu_out_4_port, alu_out(3) => 
                           alu_out_3_port, alu_out(2) => alu_out_2_port, 
                           alu_out(1) => alu_out_1_port, alu_out(0) => 
                           alu_out_0_port, alu_fw_out(31) => n_1213, 
                           alu_fw_out(30) => n_1214, alu_fw_out(29) => n_1215, 
                           alu_fw_out(28) => n_1216, alu_fw_out(27) => n_1217, 
                           alu_fw_out(26) => n_1218, alu_fw_out(25) => n_1219, 
                           alu_fw_out(24) => n_1220, alu_fw_out(23) => n_1221, 
                           alu_fw_out(22) => n_1222, alu_fw_out(21) => n_1223, 
                           alu_fw_out(20) => n_1224, alu_fw_out(19) => n_1225, 
                           alu_fw_out(18) => n_1226, alu_fw_out(17) => n_1227, 
                           alu_fw_out(16) => n_1228, alu_fw_out(15) => n_1229, 
                           alu_fw_out(14) => n_1230, alu_fw_out(13) => n_1231, 
                           alu_fw_out(12) => n_1232, alu_fw_out(11) => n_1233, 
                           alu_fw_out(10) => n_1234, alu_fw_out(9) => n_1235, 
                           alu_fw_out(8) => n_1236, alu_fw_out(7) => n_1237, 
                           alu_fw_out(6) => n_1238, alu_fw_out(5) => n_1239, 
                           alu_fw_out(4) => n_1240, alu_fw_out(3) => n_1241, 
                           alu_fw_out(2) => n_1242, alu_fw_out(1) => n_1243, 
                           alu_fw_out(0) => n_1244, r2_out(31) => 
                           aluR2_to_mem_31_port, r2_out(30) => 
                           aluR2_to_mem_30_port, r2_out(29) => 
                           aluR2_to_mem_29_port, r2_out(28) => 
                           aluR2_to_mem_28_port, r2_out(27) => 
                           aluR2_to_mem_27_port, r2_out(26) => 
                           aluR2_to_mem_26_port, r2_out(25) => 
                           aluR2_to_mem_25_port, r2_out(24) => 
                           aluR2_to_mem_24_port, r2_out(23) => 
                           aluR2_to_mem_23_port, r2_out(22) => 
                           aluR2_to_mem_22_port, r2_out(21) => 
                           aluR2_to_mem_21_port, r2_out(20) => 
                           aluR2_to_mem_20_port, r2_out(19) => 
                           aluR2_to_mem_19_port, r2_out(18) => 
                           aluR2_to_mem_18_port, r2_out(17) => 
                           aluR2_to_mem_17_port, r2_out(16) => 
                           aluR2_to_mem_16_port, r2_out(15) => 
                           aluR2_to_mem_15_port, r2_out(14) => 
                           aluR2_to_mem_14_port, r2_out(13) => 
                           aluR2_to_mem_13_port, r2_out(12) => 
                           aluR2_to_mem_12_port, r2_out(11) => 
                           aluR2_to_mem_11_port, r2_out(10) => 
                           aluR2_to_mem_10_port, r2_out(9) => 
                           aluR2_to_mem_9_port, r2_out(8) => 
                           aluR2_to_mem_8_port, r2_out(7) => 
                           aluR2_to_mem_7_port, r2_out(6) => 
                           aluR2_to_mem_6_port, r2_out(5) => 
                           aluR2_to_mem_5_port, r2_out(4) => 
                           aluR2_to_mem_4_port, r2_out(3) => 
                           aluR2_to_mem_3_port, r2_out(2) => 
                           aluR2_to_mem_2_port, r2_out(1) => 
                           aluR2_to_mem_1_port, r2_out(0) => 
                           aluR2_to_mem_0_port, b_lab_out(31) => 
                           b_from_ex_to_mem_31_port, b_lab_out(30) => 
                           b_from_ex_to_mem_30_port, b_lab_out(29) => 
                           b_from_ex_to_mem_29_port, b_lab_out(28) => 
                           b_from_ex_to_mem_28_port, b_lab_out(27) => 
                           b_from_ex_to_mem_27_port, b_lab_out(26) => 
                           b_from_ex_to_mem_26_port, b_lab_out(25) => 
                           b_from_ex_to_mem_25_port, b_lab_out(24) => 
                           b_from_ex_to_mem_24_port, b_lab_out(23) => 
                           b_from_ex_to_mem_23_port, b_lab_out(22) => 
                           b_from_ex_to_mem_22_port, b_lab_out(21) => 
                           b_from_ex_to_mem_21_port, b_lab_out(20) => 
                           b_from_ex_to_mem_20_port, b_lab_out(19) => 
                           b_from_ex_to_mem_19_port, b_lab_out(18) => 
                           b_from_ex_to_mem_18_port, b_lab_out(17) => 
                           b_from_ex_to_mem_17_port, b_lab_out(16) => 
                           b_from_ex_to_mem_16_port, b_lab_out(15) => 
                           b_from_ex_to_mem_15_port, b_lab_out(14) => 
                           b_from_ex_to_mem_14_port, b_lab_out(13) => 
                           b_from_ex_to_mem_13_port, b_lab_out(12) => 
                           b_from_ex_to_mem_12_port, b_lab_out(11) => 
                           b_from_ex_to_mem_11_port, b_lab_out(10) => 
                           b_from_ex_to_mem_10_port, b_lab_out(9) => 
                           b_from_ex_to_mem_9_port, b_lab_out(8) => 
                           b_from_ex_to_mem_8_port, b_lab_out(7) => 
                           b_from_ex_to_mem_7_port, b_lab_out(6) => 
                           b_from_ex_to_mem_6_port, b_lab_out(5) => 
                           b_from_ex_to_mem_5_port, b_lab_out(4) => 
                           b_from_ex_to_mem_4_port, b_lab_out(3) => 
                           b_from_ex_to_mem_3_port, b_lab_out(2) => 
                           b_from_ex_to_mem_2_port, b_lab_out(1) => 
                           b_from_ex_to_mem_1_port, b_lab_out(0) => 
                           b_from_ex_to_mem_0_port, pc_exe_out(31) => 
                           pc_from_ex_to_mem_31_port, pc_exe_out(30) => 
                           pc_from_ex_to_mem_30_port, pc_exe_out(29) => 
                           pc_from_ex_to_mem_29_port, pc_exe_out(28) => 
                           pc_from_ex_to_mem_28_port, pc_exe_out(27) => 
                           pc_from_ex_to_mem_27_port, pc_exe_out(26) => 
                           pc_from_ex_to_mem_26_port, pc_exe_out(25) => 
                           pc_from_ex_to_mem_25_port, pc_exe_out(24) => 
                           pc_from_ex_to_mem_24_port, pc_exe_out(23) => 
                           pc_from_ex_to_mem_23_port, pc_exe_out(22) => 
                           pc_from_ex_to_mem_22_port, pc_exe_out(21) => 
                           pc_from_ex_to_mem_21_port, pc_exe_out(20) => 
                           pc_from_ex_to_mem_20_port, pc_exe_out(19) => 
                           pc_from_ex_to_mem_19_port, pc_exe_out(18) => 
                           pc_from_ex_to_mem_18_port, pc_exe_out(17) => 
                           pc_from_ex_to_mem_17_port, pc_exe_out(16) => 
                           pc_from_ex_to_mem_16_port, pc_exe_out(15) => 
                           pc_from_ex_to_mem_15_port, pc_exe_out(14) => 
                           pc_from_ex_to_mem_14_port, pc_exe_out(13) => 
                           pc_from_ex_to_mem_13_port, pc_exe_out(12) => 
                           pc_from_ex_to_mem_12_port, pc_exe_out(11) => 
                           pc_from_ex_to_mem_11_port, pc_exe_out(10) => 
                           pc_from_ex_to_mem_10_port, pc_exe_out(9) => 
                           pc_from_ex_to_mem_9_port, pc_exe_out(8) => 
                           pc_from_ex_to_mem_8_port, pc_exe_out(7) => 
                           pc_from_ex_to_mem_7_port, pc_exe_out(6) => 
                           pc_from_ex_to_mem_6_port, pc_exe_out(5) => 
                           pc_from_ex_to_mem_5_port, pc_exe_out(4) => 
                           pc_from_ex_to_mem_4_port, pc_exe_out(3) => 
                           pc_from_ex_to_mem_3_port, pc_exe_out(2) => 
                           pc_from_ex_to_mem_2_port, pc_exe_out(1) => 
                           pc_from_ex_to_mem_1_port, pc_exe_out(0) => 
                           pc_from_ex_to_mem_0_port, rw_exe(31) => 
                           rw_from_ex_to_mem_31_port, rw_exe(30) => 
                           rw_from_ex_to_mem_30_port, rw_exe(29) => 
                           rw_from_ex_to_mem_29_port, rw_exe(28) => 
                           rw_from_ex_to_mem_28_port, rw_exe(27) => 
                           rw_from_ex_to_mem_27_port, rw_exe(26) => 
                           rw_from_ex_to_mem_26_port, rw_exe(25) => 
                           rw_from_ex_to_mem_25_port, rw_exe(24) => 
                           rw_from_ex_to_mem_24_port, rw_exe(23) => 
                           rw_from_ex_to_mem_23_port, rw_exe(22) => 
                           rw_from_ex_to_mem_22_port, rw_exe(21) => 
                           rw_from_ex_to_mem_21_port, rw_exe(20) => 
                           rw_from_ex_to_mem_20_port, rw_exe(19) => 
                           rw_from_ex_to_mem_19_port, rw_exe(18) => 
                           rw_from_ex_to_mem_18_port, rw_exe(17) => 
                           rw_from_ex_to_mem_17_port, rw_exe(16) => 
                           rw_from_ex_to_mem_16_port, rw_exe(15) => 
                           rw_from_ex_to_mem_15_port, rw_exe(14) => 
                           rw_from_ex_to_mem_14_port, rw_exe(13) => 
                           rw_from_ex_to_mem_13_port, rw_exe(12) => 
                           rw_from_ex_to_mem_12_port, rw_exe(11) => 
                           rw_from_ex_to_mem_11_port, rw_exe(10) => 
                           rw_from_ex_to_mem_10_port, rw_exe(9) => 
                           rw_from_ex_to_mem_9_port, rw_exe(8) => 
                           rw_from_ex_to_mem_8_port, rw_exe(7) => 
                           rw_from_ex_to_mem_7_port, rw_exe(6) => 
                           rw_from_ex_to_mem_6_port, rw_exe(5) => 
                           rw_from_ex_to_mem_5_port, rw_exe(4) => 
                           rw_from_ex_to_mem_4_port, rw_exe(3) => 
                           rw_from_ex_to_mem_3_port, rw_exe(2) => 
                           rw_from_ex_to_mem_2_port, rw_exe(1) => 
                           rw_from_ex_to_mem_1_port, rw_exe(0) => 
                           rw_from_ex_to_mem_0_port, j_lab_out(31) => 
                           j_from_ex_to_mem_31_port, j_lab_out(30) => 
                           j_from_ex_to_mem_30_port, j_lab_out(29) => 
                           j_from_ex_to_mem_29_port, j_lab_out(28) => 
                           j_from_ex_to_mem_28_port, j_lab_out(27) => 
                           j_from_ex_to_mem_27_port, j_lab_out(26) => 
                           j_from_ex_to_mem_26_port, j_lab_out(25) => 
                           j_from_ex_to_mem_25_port, j_lab_out(24) => 
                           j_from_ex_to_mem_24_port, j_lab_out(23) => 
                           j_from_ex_to_mem_23_port, j_lab_out(22) => 
                           j_from_ex_to_mem_22_port, j_lab_out(21) => 
                           j_from_ex_to_mem_21_port, j_lab_out(20) => 
                           j_from_ex_to_mem_20_port, j_lab_out(19) => 
                           j_from_ex_to_mem_19_port, j_lab_out(18) => 
                           j_from_ex_to_mem_18_port, j_lab_out(17) => 
                           j_from_ex_to_mem_17_port, j_lab_out(16) => 
                           j_from_ex_to_mem_16_port, j_lab_out(15) => 
                           j_from_ex_to_mem_15_port, j_lab_out(14) => 
                           j_from_ex_to_mem_14_port, j_lab_out(13) => 
                           j_from_ex_to_mem_13_port, j_lab_out(12) => 
                           j_from_ex_to_mem_12_port, j_lab_out(11) => 
                           j_from_ex_to_mem_11_port, j_lab_out(10) => 
                           j_from_ex_to_mem_10_port, j_lab_out(9) => 
                           j_from_ex_to_mem_9_port, j_lab_out(8) => 
                           j_from_ex_to_mem_8_port, j_lab_out(7) => 
                           j_from_ex_to_mem_7_port, j_lab_out(6) => 
                           j_from_ex_to_mem_6_port, j_lab_out(5) => 
                           j_from_ex_to_mem_5_port, j_lab_out(4) => 
                           j_from_ex_to_mem_4_port, j_lab_out(3) => 
                           j_from_ex_to_mem_3_port, j_lab_out(2) => 
                           j_from_ex_to_mem_2_port, j_lab_out(1) => 
                           j_from_ex_to_mem_1_port, j_lab_out(0) => 
                           j_from_ex_to_mem_0_port);
   MMU : memoryUnit_nbit32 port map( rst => n1, clk => Clk, en_reg => 
                           en_reg_mem, b_op => b_op_mem, j_op => j_op_mem, 
                           jal_op => jal_op_mem, alu_out(31) => alu_out_31_port
                           , alu_out(30) => alu_out_30_port, alu_out(29) => 
                           alu_out_29_port, alu_out(28) => alu_out_28_port, 
                           alu_out(27) => alu_out_27_port, alu_out(26) => 
                           alu_out_26_port, alu_out(25) => alu_out_25_port, 
                           alu_out(24) => alu_out_24_port, alu_out(23) => 
                           alu_out_23_port, alu_out(22) => alu_out_22_port, 
                           alu_out(21) => alu_out_21_port, alu_out(20) => 
                           alu_out_20_port, alu_out(19) => alu_out_19_port, 
                           alu_out(18) => alu_out_18_port, alu_out(17) => 
                           alu_out_17_port, alu_out(16) => alu_out_16_port, 
                           alu_out(15) => alu_out_15_port, alu_out(14) => 
                           alu_out_14_port, alu_out(13) => alu_out_13_port, 
                           alu_out(12) => alu_out_12_port, alu_out(11) => 
                           alu_out_11_port, alu_out(10) => alu_out_10_port, 
                           alu_out(9) => alu_out_9_port, alu_out(8) => 
                           alu_out_8_port, alu_out(7) => alu_out_7_port, 
                           alu_out(6) => alu_out_6_port, alu_out(5) => 
                           alu_out_5_port, alu_out(4) => alu_out_4_port, 
                           alu_out(3) => alu_out_3_port, alu_out(2) => 
                           alu_out_2_port, alu_out(1) => alu_out_1_port, 
                           alu_out(0) => alu_out_0_port, r2_out(31) => 
                           aluR2_to_mem_31_port, r2_out(30) => 
                           aluR2_to_mem_30_port, r2_out(29) => 
                           aluR2_to_mem_29_port, r2_out(28) => 
                           aluR2_to_mem_28_port, r2_out(27) => 
                           aluR2_to_mem_27_port, r2_out(26) => 
                           aluR2_to_mem_26_port, r2_out(25) => 
                           aluR2_to_mem_25_port, r2_out(24) => 
                           aluR2_to_mem_24_port, r2_out(23) => 
                           aluR2_to_mem_23_port, r2_out(22) => 
                           aluR2_to_mem_22_port, r2_out(21) => 
                           aluR2_to_mem_21_port, r2_out(20) => 
                           aluR2_to_mem_20_port, r2_out(19) => 
                           aluR2_to_mem_19_port, r2_out(18) => 
                           aluR2_to_mem_18_port, r2_out(17) => 
                           aluR2_to_mem_17_port, r2_out(16) => 
                           aluR2_to_mem_16_port, r2_out(15) => 
                           aluR2_to_mem_15_port, r2_out(14) => 
                           aluR2_to_mem_14_port, r2_out(13) => 
                           aluR2_to_mem_13_port, r2_out(12) => 
                           aluR2_to_mem_12_port, r2_out(11) => 
                           aluR2_to_mem_11_port, r2_out(10) => 
                           aluR2_to_mem_10_port, r2_out(9) => 
                           aluR2_to_mem_9_port, r2_out(8) => 
                           aluR2_to_mem_8_port, r2_out(7) => 
                           aluR2_to_mem_7_port, r2_out(6) => 
                           aluR2_to_mem_6_port, r2_out(5) => 
                           aluR2_to_mem_5_port, r2_out(4) => 
                           aluR2_to_mem_4_port, r2_out(3) => 
                           aluR2_to_mem_3_port, r2_out(2) => 
                           aluR2_to_mem_2_port, r2_out(1) => 
                           aluR2_to_mem_1_port, r2_out(0) => 
                           aluR2_to_mem_0_port, PC(31) => 
                           pc_from_ex_to_mem_31_port, PC(30) => 
                           pc_from_ex_to_mem_30_port, PC(29) => 
                           pc_from_ex_to_mem_29_port, PC(28) => 
                           pc_from_ex_to_mem_28_port, PC(27) => 
                           pc_from_ex_to_mem_27_port, PC(26) => 
                           pc_from_ex_to_mem_26_port, PC(25) => 
                           pc_from_ex_to_mem_25_port, PC(24) => 
                           pc_from_ex_to_mem_24_port, PC(23) => 
                           pc_from_ex_to_mem_23_port, PC(22) => 
                           pc_from_ex_to_mem_22_port, PC(21) => 
                           pc_from_ex_to_mem_21_port, PC(20) => 
                           pc_from_ex_to_mem_20_port, PC(19) => 
                           pc_from_ex_to_mem_19_port, PC(18) => 
                           pc_from_ex_to_mem_18_port, PC(17) => 
                           pc_from_ex_to_mem_17_port, PC(16) => 
                           pc_from_ex_to_mem_16_port, PC(15) => 
                           pc_from_ex_to_mem_15_port, PC(14) => 
                           pc_from_ex_to_mem_14_port, PC(13) => 
                           pc_from_ex_to_mem_13_port, PC(12) => 
                           pc_from_ex_to_mem_12_port, PC(11) => 
                           pc_from_ex_to_mem_11_port, PC(10) => 
                           pc_from_ex_to_mem_10_port, PC(9) => 
                           pc_from_ex_to_mem_9_port, PC(8) => 
                           pc_from_ex_to_mem_8_port, PC(7) => 
                           pc_from_ex_to_mem_7_port, PC(6) => 
                           pc_from_ex_to_mem_6_port, PC(5) => 
                           pc_from_ex_to_mem_5_port, PC(4) => 
                           pc_from_ex_to_mem_4_port, PC(3) => 
                           pc_from_ex_to_mem_3_port, PC(2) => 
                           pc_from_ex_to_mem_2_port, PC(1) => 
                           pc_from_ex_to_mem_1_port, PC(0) => 
                           pc_from_ex_to_mem_0_port, lab_b(31) => 
                           b_from_ex_to_mem_31_port, lab_b(30) => 
                           b_from_ex_to_mem_30_port, lab_b(29) => 
                           b_from_ex_to_mem_29_port, lab_b(28) => 
                           b_from_ex_to_mem_28_port, lab_b(27) => 
                           b_from_ex_to_mem_27_port, lab_b(26) => 
                           b_from_ex_to_mem_26_port, lab_b(25) => 
                           b_from_ex_to_mem_25_port, lab_b(24) => 
                           b_from_ex_to_mem_24_port, lab_b(23) => 
                           b_from_ex_to_mem_23_port, lab_b(22) => 
                           b_from_ex_to_mem_22_port, lab_b(21) => 
                           b_from_ex_to_mem_21_port, lab_b(20) => 
                           b_from_ex_to_mem_20_port, lab_b(19) => 
                           b_from_ex_to_mem_19_port, lab_b(18) => 
                           b_from_ex_to_mem_18_port, lab_b(17) => 
                           b_from_ex_to_mem_17_port, lab_b(16) => 
                           b_from_ex_to_mem_16_port, lab_b(15) => 
                           b_from_ex_to_mem_15_port, lab_b(14) => 
                           b_from_ex_to_mem_14_port, lab_b(13) => 
                           b_from_ex_to_mem_13_port, lab_b(12) => 
                           b_from_ex_to_mem_12_port, lab_b(11) => 
                           b_from_ex_to_mem_11_port, lab_b(10) => 
                           b_from_ex_to_mem_10_port, lab_b(9) => 
                           b_from_ex_to_mem_9_port, lab_b(8) => 
                           b_from_ex_to_mem_8_port, lab_b(7) => 
                           b_from_ex_to_mem_7_port, lab_b(6) => 
                           b_from_ex_to_mem_6_port, lab_b(5) => 
                           b_from_ex_to_mem_5_port, lab_b(4) => 
                           b_from_ex_to_mem_4_port, lab_b(3) => 
                           b_from_ex_to_mem_3_port, lab_b(2) => 
                           b_from_ex_to_mem_2_port, lab_b(1) => 
                           b_from_ex_to_mem_1_port, lab_b(0) => 
                           b_from_ex_to_mem_0_port, lab_j(31) => 
                           j_from_ex_to_mem_31_port, lab_j(30) => 
                           j_from_ex_to_mem_30_port, lab_j(29) => 
                           j_from_ex_to_mem_29_port, lab_j(28) => 
                           j_from_ex_to_mem_28_port, lab_j(27) => 
                           j_from_ex_to_mem_27_port, lab_j(26) => 
                           j_from_ex_to_mem_26_port, lab_j(25) => 
                           j_from_ex_to_mem_25_port, lab_j(24) => 
                           j_from_ex_to_mem_24_port, lab_j(23) => 
                           j_from_ex_to_mem_23_port, lab_j(22) => 
                           j_from_ex_to_mem_22_port, lab_j(21) => 
                           j_from_ex_to_mem_21_port, lab_j(20) => 
                           j_from_ex_to_mem_20_port, lab_j(19) => 
                           j_from_ex_to_mem_19_port, lab_j(18) => 
                           j_from_ex_to_mem_18_port, lab_j(17) => 
                           j_from_ex_to_mem_17_port, lab_j(16) => 
                           j_from_ex_to_mem_16_port, lab_j(15) => 
                           j_from_ex_to_mem_15_port, lab_j(14) => 
                           j_from_ex_to_mem_14_port, lab_j(13) => 
                           j_from_ex_to_mem_13_port, lab_j(12) => 
                           j_from_ex_to_mem_12_port, lab_j(11) => 
                           j_from_ex_to_mem_11_port, lab_j(10) => 
                           j_from_ex_to_mem_10_port, lab_j(9) => 
                           j_from_ex_to_mem_9_port, lab_j(8) => 
                           j_from_ex_to_mem_8_port, lab_j(7) => 
                           j_from_ex_to_mem_7_port, lab_j(6) => 
                           j_from_ex_to_mem_6_port, lab_j(5) => 
                           j_from_ex_to_mem_5_port, lab_j(4) => 
                           j_from_ex_to_mem_4_port, lab_j(3) => 
                           j_from_ex_to_mem_3_port, lab_j(2) => 
                           j_from_ex_to_mem_2_port, lab_j(1) => 
                           j_from_ex_to_mem_1_port, lab_j(0) => 
                           j_from_ex_to_mem_0_port, rw_exe(31) => 
                           rw_from_ex_to_mem_31_port, rw_exe(30) => 
                           rw_from_ex_to_mem_30_port, rw_exe(29) => 
                           rw_from_ex_to_mem_29_port, rw_exe(28) => 
                           rw_from_ex_to_mem_28_port, rw_exe(27) => 
                           rw_from_ex_to_mem_27_port, rw_exe(26) => 
                           rw_from_ex_to_mem_26_port, rw_exe(25) => 
                           rw_from_ex_to_mem_25_port, rw_exe(24) => 
                           rw_from_ex_to_mem_24_port, rw_exe(23) => 
                           rw_from_ex_to_mem_23_port, rw_exe(22) => 
                           rw_from_ex_to_mem_22_port, rw_exe(21) => 
                           rw_from_ex_to_mem_21_port, rw_exe(20) => 
                           rw_from_ex_to_mem_20_port, rw_exe(19) => 
                           rw_from_ex_to_mem_19_port, rw_exe(18) => 
                           rw_from_ex_to_mem_18_port, rw_exe(17) => 
                           rw_from_ex_to_mem_17_port, rw_exe(16) => 
                           rw_from_ex_to_mem_16_port, rw_exe(15) => 
                           rw_from_ex_to_mem_15_port, rw_exe(14) => 
                           rw_from_ex_to_mem_14_port, rw_exe(13) => 
                           rw_from_ex_to_mem_13_port, rw_exe(12) => 
                           rw_from_ex_to_mem_12_port, rw_exe(11) => 
                           rw_from_ex_to_mem_11_port, rw_exe(10) => 
                           rw_from_ex_to_mem_10_port, rw_exe(9) => 
                           rw_from_ex_to_mem_9_port, rw_exe(8) => 
                           rw_from_ex_to_mem_8_port, rw_exe(7) => 
                           rw_from_ex_to_mem_7_port, rw_exe(6) => 
                           rw_from_ex_to_mem_6_port, rw_exe(5) => 
                           rw_from_ex_to_mem_5_port, rw_exe(4) => 
                           rw_from_ex_to_mem_4_port, rw_exe(3) => 
                           rw_from_ex_to_mem_3_port, rw_exe(2) => 
                           rw_from_ex_to_mem_2_port, rw_exe(1) => 
                           rw_from_ex_to_mem_1_port, rw_exe(0) => 
                           rw_from_ex_to_mem_0_port, dataout_from_mem(31) => 
                           dataout_from_mem(31), dataout_from_mem(30) => 
                           dataout_from_mem(30), dataout_from_mem(29) => 
                           dataout_from_mem(29), dataout_from_mem(28) => 
                           dataout_from_mem(28), dataout_from_mem(27) => 
                           dataout_from_mem(27), dataout_from_mem(26) => 
                           dataout_from_mem(26), dataout_from_mem(25) => 
                           dataout_from_mem(25), dataout_from_mem(24) => 
                           dataout_from_mem(24), dataout_from_mem(23) => 
                           dataout_from_mem(23), dataout_from_mem(22) => 
                           dataout_from_mem(22), dataout_from_mem(21) => 
                           dataout_from_mem(21), dataout_from_mem(20) => 
                           dataout_from_mem(20), dataout_from_mem(19) => 
                           dataout_from_mem(19), dataout_from_mem(18) => 
                           dataout_from_mem(18), dataout_from_mem(17) => 
                           dataout_from_mem(17), dataout_from_mem(16) => 
                           dataout_from_mem(16), dataout_from_mem(15) => 
                           dataout_from_mem(15), dataout_from_mem(14) => 
                           dataout_from_mem(14), dataout_from_mem(13) => 
                           dataout_from_mem(13), dataout_from_mem(12) => 
                           dataout_from_mem(12), dataout_from_mem(11) => 
                           dataout_from_mem(11), dataout_from_mem(10) => 
                           dataout_from_mem(10), dataout_from_mem(9) => 
                           dataout_from_mem(9), dataout_from_mem(8) => 
                           dataout_from_mem(8), dataout_from_mem(7) => 
                           dataout_from_mem(7), dataout_from_mem(6) => 
                           dataout_from_mem(6), dataout_from_mem(5) => 
                           dataout_from_mem(5), dataout_from_mem(4) => 
                           dataout_from_mem(4), dataout_from_mem(3) => 
                           dataout_from_mem(3), dataout_from_mem(2) => 
                           dataout_from_mem(2), dataout_from_mem(1) => 
                           dataout_from_mem(1), dataout_from_mem(0) => 
                           dataout_from_mem(0), addr_mem(31) => addr_mem(31), 
                           addr_mem(30) => addr_mem(30), addr_mem(29) => 
                           addr_mem(29), addr_mem(28) => addr_mem(28), 
                           addr_mem(27) => addr_mem(27), addr_mem(26) => 
                           addr_mem(26), addr_mem(25) => addr_mem(25), 
                           addr_mem(24) => addr_mem(24), addr_mem(23) => 
                           addr_mem(23), addr_mem(22) => addr_mem(22), 
                           addr_mem(21) => addr_mem(21), addr_mem(20) => 
                           addr_mem(20), addr_mem(19) => addr_mem(19), 
                           addr_mem(18) => addr_mem(18), addr_mem(17) => 
                           addr_mem(17), addr_mem(16) => addr_mem(16), 
                           addr_mem(15) => addr_mem(15), addr_mem(14) => 
                           addr_mem(14), addr_mem(13) => addr_mem(13), 
                           addr_mem(12) => addr_mem(12), addr_mem(11) => 
                           addr_mem(11), addr_mem(10) => addr_mem(10), 
                           addr_mem(9) => addr_mem(9), addr_mem(8) => 
                           addr_mem(8), addr_mem(7) => addr_mem(7), addr_mem(6)
                           => addr_mem(6), addr_mem(5) => addr_mem(5), 
                           addr_mem(4) => addr_mem(4), addr_mem(3) => 
                           addr_mem(3), addr_mem(2) => addr_mem(2), addr_mem(1)
                           => addr_mem(1), addr_mem(0) => addr_mem(0), 
                           datain_mem(31) => datain_mem(31), datain_mem(30) => 
                           datain_mem(30), datain_mem(29) => datain_mem(29), 
                           datain_mem(28) => datain_mem(28), datain_mem(27) => 
                           datain_mem(27), datain_mem(26) => datain_mem(26), 
                           datain_mem(25) => datain_mem(25), datain_mem(24) => 
                           datain_mem(24), datain_mem(23) => datain_mem(23), 
                           datain_mem(22) => datain_mem(22), datain_mem(21) => 
                           datain_mem(21), datain_mem(20) => datain_mem(20), 
                           datain_mem(19) => datain_mem(19), datain_mem(18) => 
                           datain_mem(18), datain_mem(17) => datain_mem(17), 
                           datain_mem(16) => datain_mem(16), datain_mem(15) => 
                           datain_mem(15), datain_mem(14) => datain_mem(14), 
                           datain_mem(13) => datain_mem(13), datain_mem(12) => 
                           datain_mem(12), datain_mem(11) => datain_mem(11), 
                           datain_mem(10) => datain_mem(10), datain_mem(9) => 
                           datain_mem(9), datain_mem(8) => datain_mem(8), 
                           datain_mem(7) => datain_mem(7), datain_mem(6) => 
                           datain_mem(6), datain_mem(5) => datain_mem(5), 
                           datain_mem(4) => datain_mem(4), datain_mem(3) => 
                           datain_mem(3), datain_mem(2) => datain_mem(2), 
                           datain_mem(1) => datain_mem(1), datain_mem(0) => 
                           datain_mem(0), next_PC(31) => 
                           pc_from_mem_to_fetch_31_port, next_PC(30) => 
                           pc_from_mem_to_fetch_30_port, next_PC(29) => 
                           pc_from_mem_to_fetch_29_port, next_PC(28) => 
                           pc_from_mem_to_fetch_28_port, next_PC(27) => 
                           pc_from_mem_to_fetch_27_port, next_PC(26) => 
                           pc_from_mem_to_fetch_26_port, next_PC(25) => 
                           pc_from_mem_to_fetch_25_port, next_PC(24) => 
                           pc_from_mem_to_fetch_24_port, next_PC(23) => 
                           pc_from_mem_to_fetch_23_port, next_PC(22) => 
                           pc_from_mem_to_fetch_22_port, next_PC(21) => 
                           pc_from_mem_to_fetch_21_port, next_PC(20) => 
                           pc_from_mem_to_fetch_20_port, next_PC(19) => 
                           pc_from_mem_to_fetch_19_port, next_PC(18) => 
                           pc_from_mem_to_fetch_18_port, next_PC(17) => 
                           pc_from_mem_to_fetch_17_port, next_PC(16) => 
                           pc_from_mem_to_fetch_16_port, next_PC(15) => 
                           pc_from_mem_to_fetch_15_port, next_PC(14) => 
                           pc_from_mem_to_fetch_14_port, next_PC(13) => 
                           pc_from_mem_to_fetch_13_port, next_PC(12) => 
                           pc_from_mem_to_fetch_12_port, next_PC(11) => 
                           pc_from_mem_to_fetch_11_port, next_PC(10) => 
                           pc_from_mem_to_fetch_10_port, next_PC(9) => 
                           pc_from_mem_to_fetch_9_port, next_PC(8) => 
                           pc_from_mem_to_fetch_8_port, next_PC(7) => 
                           pc_from_mem_to_fetch_7_port, next_PC(6) => 
                           pc_from_mem_to_fetch_6_port, next_PC(5) => 
                           pc_from_mem_to_fetch_5_port, next_PC(4) => 
                           pc_from_mem_to_fetch_4_port, next_PC(3) => 
                           pc_from_mem_to_fetch_3_port, next_PC(2) => 
                           pc_from_mem_to_fetch_2_port, next_PC(1) => 
                           pc_from_mem_to_fetch_1_port, next_PC(0) => 
                           pc_from_mem_to_fetch_0_port, alu_out_mem(31) => 
                           alu_out_mem_31_port, alu_out_mem(30) => 
                           alu_out_mem_30_port, alu_out_mem(29) => 
                           alu_out_mem_29_port, alu_out_mem(28) => 
                           alu_out_mem_28_port, alu_out_mem(27) => 
                           alu_out_mem_27_port, alu_out_mem(26) => 
                           alu_out_mem_26_port, alu_out_mem(25) => 
                           alu_out_mem_25_port, alu_out_mem(24) => 
                           alu_out_mem_24_port, alu_out_mem(23) => 
                           alu_out_mem_23_port, alu_out_mem(22) => 
                           alu_out_mem_22_port, alu_out_mem(21) => 
                           alu_out_mem_21_port, alu_out_mem(20) => 
                           alu_out_mem_20_port, alu_out_mem(19) => 
                           alu_out_mem_19_port, alu_out_mem(18) => 
                           alu_out_mem_18_port, alu_out_mem(17) => 
                           alu_out_mem_17_port, alu_out_mem(16) => 
                           alu_out_mem_16_port, alu_out_mem(15) => 
                           alu_out_mem_15_port, alu_out_mem(14) => 
                           alu_out_mem_14_port, alu_out_mem(13) => 
                           alu_out_mem_13_port, alu_out_mem(12) => 
                           alu_out_mem_12_port, alu_out_mem(11) => 
                           alu_out_mem_11_port, alu_out_mem(10) => 
                           alu_out_mem_10_port, alu_out_mem(9) => 
                           alu_out_mem_9_port, alu_out_mem(8) => 
                           alu_out_mem_8_port, alu_out_mem(7) => 
                           alu_out_mem_7_port, alu_out_mem(6) => 
                           alu_out_mem_6_port, alu_out_mem(5) => 
                           alu_out_mem_5_port, alu_out_mem(4) => 
                           alu_out_mem_4_port, alu_out_mem(3) => 
                           alu_out_mem_3_port, alu_out_mem(2) => 
                           alu_out_mem_2_port, alu_out_mem(1) => 
                           alu_out_mem_1_port, alu_out_mem(0) => 
                           alu_out_mem_0_port, rw_mem(31) => n_1245, rw_mem(30)
                           => n_1246, rw_mem(29) => n_1247, rw_mem(28) => 
                           n_1248, rw_mem(27) => n_1249, rw_mem(26) => n_1250, 
                           rw_mem(25) => n_1251, rw_mem(24) => n_1252, 
                           rw_mem(23) => n_1253, rw_mem(22) => n_1254, 
                           rw_mem(21) => n_1255, rw_mem(20) => n_1256, 
                           rw_mem(19) => n_1257, rw_mem(18) => n_1258, 
                           rw_mem(17) => n_1259, rw_mem(16) => n_1260, 
                           rw_mem(15) => n_1261, rw_mem(14) => n_1262, 
                           rw_mem(13) => n_1263, rw_mem(12) => n_1264, 
                           rw_mem(11) => n_1265, rw_mem(10) => n_1266, 
                           rw_mem(9) => n_1267, rw_mem(8) => n_1268, rw_mem(7) 
                           => n_1269, rw_mem(6) => n_1270, rw_mem(5) => n_1271,
                           rw_mem(4) => ADD_RW_4_port, rw_mem(3) => 
                           ADD_RW_3_port, rw_mem(2) => ADD_RW_2_port, rw_mem(1)
                           => ADD_RW_1_port, rw_mem(0) => ADD_RW_0_port, 
                           data_out(31) => data_from_mem_to_wb_31_port, 
                           data_out(30) => data_from_mem_to_wb_30_port, 
                           data_out(29) => data_from_mem_to_wb_29_port, 
                           data_out(28) => data_from_mem_to_wb_28_port, 
                           data_out(27) => data_from_mem_to_wb_27_port, 
                           data_out(26) => data_from_mem_to_wb_26_port, 
                           data_out(25) => data_from_mem_to_wb_25_port, 
                           data_out(24) => data_from_mem_to_wb_24_port, 
                           data_out(23) => data_from_mem_to_wb_23_port, 
                           data_out(22) => data_from_mem_to_wb_22_port, 
                           data_out(21) => data_from_mem_to_wb_21_port, 
                           data_out(20) => data_from_mem_to_wb_20_port, 
                           data_out(19) => data_from_mem_to_wb_19_port, 
                           data_out(18) => data_from_mem_to_wb_18_port, 
                           data_out(17) => data_from_mem_to_wb_17_port, 
                           data_out(16) => data_from_mem_to_wb_16_port, 
                           data_out(15) => data_from_mem_to_wb_15_port, 
                           data_out(14) => data_from_mem_to_wb_14_port, 
                           data_out(13) => data_from_mem_to_wb_13_port, 
                           data_out(12) => data_from_mem_to_wb_12_port, 
                           data_out(11) => data_from_mem_to_wb_11_port, 
                           data_out(10) => data_from_mem_to_wb_10_port, 
                           data_out(9) => data_from_mem_to_wb_9_port, 
                           data_out(8) => data_from_mem_to_wb_8_port, 
                           data_out(7) => data_from_mem_to_wb_7_port, 
                           data_out(6) => data_from_mem_to_wb_6_port, 
                           data_out(5) => data_from_mem_to_wb_5_port, 
                           data_out(4) => data_from_mem_to_wb_4_port, 
                           data_out(3) => data_from_mem_to_wb_3_port, 
                           data_out(2) => data_from_mem_to_wb_2_port, 
                           data_out(1) => data_from_mem_to_wb_1_port, 
                           data_out(0) => data_from_mem_to_wb_0_port);
   WBU : writeBackUnit_nbit32 port map( MemtoReg => MemtoReg_wb, ReadData(31) 
                           => data_from_mem_to_wb_31_port, ReadData(30) => 
                           data_from_mem_to_wb_30_port, ReadData(29) => 
                           data_from_mem_to_wb_29_port, ReadData(28) => 
                           data_from_mem_to_wb_28_port, ReadData(27) => 
                           data_from_mem_to_wb_27_port, ReadData(26) => 
                           data_from_mem_to_wb_26_port, ReadData(25) => 
                           data_from_mem_to_wb_25_port, ReadData(24) => 
                           data_from_mem_to_wb_24_port, ReadData(23) => 
                           data_from_mem_to_wb_23_port, ReadData(22) => 
                           data_from_mem_to_wb_22_port, ReadData(21) => 
                           data_from_mem_to_wb_21_port, ReadData(20) => 
                           data_from_mem_to_wb_20_port, ReadData(19) => 
                           data_from_mem_to_wb_19_port, ReadData(18) => 
                           data_from_mem_to_wb_18_port, ReadData(17) => 
                           data_from_mem_to_wb_17_port, ReadData(16) => 
                           data_from_mem_to_wb_16_port, ReadData(15) => 
                           data_from_mem_to_wb_15_port, ReadData(14) => 
                           data_from_mem_to_wb_14_port, ReadData(13) => 
                           data_from_mem_to_wb_13_port, ReadData(12) => 
                           data_from_mem_to_wb_12_port, ReadData(11) => 
                           data_from_mem_to_wb_11_port, ReadData(10) => 
                           data_from_mem_to_wb_10_port, ReadData(9) => 
                           data_from_mem_to_wb_9_port, ReadData(8) => 
                           data_from_mem_to_wb_8_port, ReadData(7) => 
                           data_from_mem_to_wb_7_port, ReadData(6) => 
                           data_from_mem_to_wb_6_port, ReadData(5) => 
                           data_from_mem_to_wb_5_port, ReadData(4) => 
                           data_from_mem_to_wb_4_port, ReadData(3) => 
                           data_from_mem_to_wb_3_port, ReadData(2) => 
                           data_from_mem_to_wb_2_port, ReadData(1) => 
                           data_from_mem_to_wb_1_port, ReadData(0) => 
                           data_from_mem_to_wb_0_port, AluResult(31) => 
                           alu_out_mem_31_port, AluResult(30) => 
                           alu_out_mem_30_port, AluResult(29) => 
                           alu_out_mem_29_port, AluResult(28) => 
                           alu_out_mem_28_port, AluResult(27) => 
                           alu_out_mem_27_port, AluResult(26) => 
                           alu_out_mem_26_port, AluResult(25) => 
                           alu_out_mem_25_port, AluResult(24) => 
                           alu_out_mem_24_port, AluResult(23) => 
                           alu_out_mem_23_port, AluResult(22) => 
                           alu_out_mem_22_port, AluResult(21) => 
                           alu_out_mem_21_port, AluResult(20) => 
                           alu_out_mem_20_port, AluResult(19) => 
                           alu_out_mem_19_port, AluResult(18) => 
                           alu_out_mem_18_port, AluResult(17) => 
                           alu_out_mem_17_port, AluResult(16) => 
                           alu_out_mem_16_port, AluResult(15) => 
                           alu_out_mem_15_port, AluResult(14) => 
                           alu_out_mem_14_port, AluResult(13) => 
                           alu_out_mem_13_port, AluResult(12) => 
                           alu_out_mem_12_port, AluResult(11) => 
                           alu_out_mem_11_port, AluResult(10) => 
                           alu_out_mem_10_port, AluResult(9) => 
                           alu_out_mem_9_port, AluResult(8) => 
                           alu_out_mem_8_port, AluResult(7) => 
                           alu_out_mem_7_port, AluResult(6) => 
                           alu_out_mem_6_port, AluResult(5) => 
                           alu_out_mem_5_port, AluResult(4) => 
                           alu_out_mem_4_port, AluResult(3) => 
                           alu_out_mem_3_port, AluResult(2) => 
                           alu_out_mem_2_port, AluResult(1) => 
                           alu_out_mem_1_port, AluResult(0) => 
                           alu_out_mem_0_port, WriteData(31) => 
                           pipe_out_31_port, WriteData(30) => pipe_out_30_port,
                           WriteData(29) => pipe_out_29_port, WriteData(28) => 
                           pipe_out_28_port, WriteData(27) => pipe_out_27_port,
                           WriteData(26) => pipe_out_26_port, WriteData(25) => 
                           pipe_out_25_port, WriteData(24) => pipe_out_24_port,
                           WriteData(23) => pipe_out_23_port, WriteData(22) => 
                           pipe_out_22_port, WriteData(21) => pipe_out_21_port,
                           WriteData(20) => pipe_out_20_port, WriteData(19) => 
                           pipe_out_19_port, WriteData(18) => pipe_out_18_port,
                           WriteData(17) => pipe_out_17_port, WriteData(16) => 
                           pipe_out_16_port, WriteData(15) => pipe_out_15_port,
                           WriteData(14) => pipe_out_14_port, WriteData(13) => 
                           pipe_out_13_port, WriteData(12) => pipe_out_12_port,
                           WriteData(11) => pipe_out_11_port, WriteData(10) => 
                           pipe_out_10_port, WriteData(9) => pipe_out_9_port, 
                           WriteData(8) => pipe_out_8_port, WriteData(7) => 
                           pipe_out_7_port, WriteData(6) => pipe_out_6_port, 
                           WriteData(5) => pipe_out_5_port, WriteData(4) => 
                           pipe_out_4_port, WriteData(3) => pipe_out_3_port, 
                           WriteData(2) => pipe_out_2_port, WriteData(1) => 
                           pipe_out_1_port, WriteData(0) => pipe_out_0_port);
   U1 : BUF_X2 port map( A => Rst, Z => n1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_nbit32.all;

entity DLX_nbit32 is

   port( Clk, Rst : in std_logic;  dout_IRAM : in std_logic_vector (31 downto 
         0);  addr_IRAM : out std_logic_vector (31 downto 0);  MEM_EN_MEM, 
         RD_MEM, WR_MEM : out std_logic;  dataout_from_mem : in 
         std_logic_vector (31 downto 0);  addr_mem, datain_mem, dlx_data_out : 
         out std_logic_vector (31 downto 0));

end DLX_nbit32;

architecture SYN_dlx_rtl of DLX_nbit32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE45_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13
      port( Clk, Rst, En : in std_logic;  IR_opcode : in std_logic_vector (5 
            downto 0);  IR_func : in std_logic_vector (10 downto 0);  PC_OP, 
            EN_REG_IF, EN_REG_ID, RD1, RD2, SEL_EX, EN_REG_EX, SEL_MUX_RW : out
            std_logic;  ALU_OPCODE : out std_logic_vector (3 downto 0);  
            EN_REG_MEM, MEM_EN_MEM, RD_MEM, WR_MEM, B_OP_MEM, J_OP_MEM, 
            JAL_OP_MEM, MEM_TO_REG_WB, WR : out std_logic);
   end component;
   
   component flip_flop_1
      port( D, CK, Enable_n, RESET_n : in std_logic;  Q : out std_logic);
   end component;
   
   component flip_flop_0
      port( D, CK, Enable_n, RESET_n : in std_logic;  Q : out std_logic);
   end component;
   
   component datapath_nbit32
      port( Clk, Rst, PC_op, en_reg_if, RD1, RD2 : in std_logic;  dout_IRAM : 
            in std_logic_vector (31 downto 0);  addr_IRAM : out 
            std_logic_vector (31 downto 0);  en_reg_id, WR : in std_logic;  
            Opcode : out std_logic_vector (5 downto 0);  Func : out 
            std_logic_vector (10 downto 0);  sel_ex, sel_mux_rw, en_reg_ex : in
            std_logic;  alu_sel : in std_logic_vector (3 downto 0);  en_reg_mem
            : in std_logic;  dataout_from_mem : in std_logic_vector (31 downto 
            0);  addr_mem, datain_mem : out std_logic_vector (31 downto 0);  
            b_op_mem, j_op_mem, jal_op_mem, MemtoReg_wb : in std_logic;  
            pipe_out : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, PC_op_i, en_reg_if_i, RD1_i, RD2_i, 
      en_reg_id_i, WR_i, Opcode_i_5_port, Opcode_i_4_port, Opcode_i_3_port, 
      Opcode_i_2_port, Opcode_i_1_port, Opcode_i_0_port, Func_i_10_port, 
      Func_i_9_port, Func_i_8_port, Func_i_7_port, Func_i_6_port, Func_i_5_port
      , Func_i_4_port, Func_i_3_port, Func_i_2_port, Func_i_1_port, 
      Func_i_0_port, sel_ex_i, sel_mux_rw_i, en_reg_ex_i, alu_sel_i_3_port, 
      alu_sel_i_2_port, alu_sel_i_1_port, alu_sel_i_0_port, en_reg_mem_i, 
      b_op_mem_i, j_op_mem_i, jal_op_mem_i, MemtoReg_wb_i, CU_en1, CU_en2, n4, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   WR_i <= '0';
   jal_op_mem_i <= '0';
   j_op_mem_i <= '0';
   b_op_mem_i <= '0';
   WR_MEM <= '0';
   RD_MEM <= '0';
   sel_mux_rw_i <= '0';
   sel_ex_i <= '0';
   PC_op_i <= '0';
   DataPath_dlx : datapath_nbit32 port map( Clk => Clk, Rst => Rst, PC_op => 
                           PC_op_i, en_reg_if => en_reg_if_i, RD1 => RD1_i, RD2
                           => RD2_i, dout_IRAM(31) => dout_IRAM(31), 
                           dout_IRAM(30) => dout_IRAM(30), dout_IRAM(29) => 
                           dout_IRAM(29), dout_IRAM(28) => dout_IRAM(28), 
                           dout_IRAM(27) => dout_IRAM(27), dout_IRAM(26) => 
                           dout_IRAM(26), dout_IRAM(25) => dout_IRAM(25), 
                           dout_IRAM(24) => dout_IRAM(24), dout_IRAM(23) => 
                           dout_IRAM(23), dout_IRAM(22) => dout_IRAM(22), 
                           dout_IRAM(21) => dout_IRAM(21), dout_IRAM(20) => 
                           dout_IRAM(20), dout_IRAM(19) => dout_IRAM(19), 
                           dout_IRAM(18) => dout_IRAM(18), dout_IRAM(17) => 
                           dout_IRAM(17), dout_IRAM(16) => dout_IRAM(16), 
                           dout_IRAM(15) => dout_IRAM(15), dout_IRAM(14) => 
                           dout_IRAM(14), dout_IRAM(13) => dout_IRAM(13), 
                           dout_IRAM(12) => dout_IRAM(12), dout_IRAM(11) => 
                           dout_IRAM(11), dout_IRAM(10) => dout_IRAM(10), 
                           dout_IRAM(9) => dout_IRAM(9), dout_IRAM(8) => 
                           dout_IRAM(8), dout_IRAM(7) => dout_IRAM(7), 
                           dout_IRAM(6) => dout_IRAM(6), dout_IRAM(5) => 
                           dout_IRAM(5), dout_IRAM(4) => dout_IRAM(4), 
                           dout_IRAM(3) => dout_IRAM(3), dout_IRAM(2) => 
                           dout_IRAM(2), dout_IRAM(1) => dout_IRAM(1), 
                           dout_IRAM(0) => dout_IRAM(0), addr_IRAM(31) => 
                           addr_IRAM(31), addr_IRAM(30) => addr_IRAM(30), 
                           addr_IRAM(29) => addr_IRAM(29), addr_IRAM(28) => 
                           addr_IRAM(28), addr_IRAM(27) => addr_IRAM(27), 
                           addr_IRAM(26) => addr_IRAM(26), addr_IRAM(25) => 
                           addr_IRAM(25), addr_IRAM(24) => addr_IRAM(24), 
                           addr_IRAM(23) => addr_IRAM(23), addr_IRAM(22) => 
                           addr_IRAM(22), addr_IRAM(21) => addr_IRAM(21), 
                           addr_IRAM(20) => addr_IRAM(20), addr_IRAM(19) => 
                           addr_IRAM(19), addr_IRAM(18) => addr_IRAM(18), 
                           addr_IRAM(17) => addr_IRAM(17), addr_IRAM(16) => 
                           addr_IRAM(16), addr_IRAM(15) => addr_IRAM(15), 
                           addr_IRAM(14) => addr_IRAM(14), addr_IRAM(13) => 
                           addr_IRAM(13), addr_IRAM(12) => addr_IRAM(12), 
                           addr_IRAM(11) => addr_IRAM(11), addr_IRAM(10) => 
                           addr_IRAM(10), addr_IRAM(9) => addr_IRAM(9), 
                           addr_IRAM(8) => addr_IRAM(8), addr_IRAM(7) => 
                           addr_IRAM(7), addr_IRAM(6) => addr_IRAM(6), 
                           addr_IRAM(5) => addr_IRAM(5), addr_IRAM(4) => 
                           addr_IRAM(4), addr_IRAM(3) => addr_IRAM(3), 
                           addr_IRAM(2) => addr_IRAM(2), addr_IRAM(1) => 
                           addr_IRAM(1), addr_IRAM(0) => addr_IRAM(0), 
                           en_reg_id => en_reg_id_i, WR => WR_i, Opcode(5) => 
                           Opcode_i_5_port, Opcode(4) => Opcode_i_4_port, 
                           Opcode(3) => Opcode_i_3_port, Opcode(2) => 
                           Opcode_i_2_port, Opcode(1) => Opcode_i_1_port, 
                           Opcode(0) => Opcode_i_0_port, Func(10) => 
                           Func_i_10_port, Func(9) => Func_i_9_port, Func(8) =>
                           Func_i_8_port, Func(7) => Func_i_7_port, Func(6) => 
                           Func_i_6_port, Func(5) => Func_i_5_port, Func(4) => 
                           Func_i_4_port, Func(3) => Func_i_3_port, Func(2) => 
                           Func_i_2_port, Func(1) => Func_i_1_port, Func(0) => 
                           Func_i_0_port, sel_ex => sel_ex_i, sel_mux_rw => 
                           sel_mux_rw_i, en_reg_ex => en_reg_ex_i, alu_sel(3) 
                           => alu_sel_i_3_port, alu_sel(2) => alu_sel_i_2_port,
                           alu_sel(1) => alu_sel_i_1_port, alu_sel(0) => 
                           alu_sel_i_0_port, en_reg_mem => en_reg_mem_i, 
                           dataout_from_mem(31) => dataout_from_mem(31), 
                           dataout_from_mem(30) => dataout_from_mem(30), 
                           dataout_from_mem(29) => dataout_from_mem(29), 
                           dataout_from_mem(28) => dataout_from_mem(28), 
                           dataout_from_mem(27) => dataout_from_mem(27), 
                           dataout_from_mem(26) => dataout_from_mem(26), 
                           dataout_from_mem(25) => dataout_from_mem(25), 
                           dataout_from_mem(24) => dataout_from_mem(24), 
                           dataout_from_mem(23) => dataout_from_mem(23), 
                           dataout_from_mem(22) => dataout_from_mem(22), 
                           dataout_from_mem(21) => dataout_from_mem(21), 
                           dataout_from_mem(20) => dataout_from_mem(20), 
                           dataout_from_mem(19) => dataout_from_mem(19), 
                           dataout_from_mem(18) => dataout_from_mem(18), 
                           dataout_from_mem(17) => dataout_from_mem(17), 
                           dataout_from_mem(16) => dataout_from_mem(16), 
                           dataout_from_mem(15) => dataout_from_mem(15), 
                           dataout_from_mem(14) => dataout_from_mem(14), 
                           dataout_from_mem(13) => dataout_from_mem(13), 
                           dataout_from_mem(12) => dataout_from_mem(12), 
                           dataout_from_mem(11) => dataout_from_mem(11), 
                           dataout_from_mem(10) => dataout_from_mem(10), 
                           dataout_from_mem(9) => dataout_from_mem(9), 
                           dataout_from_mem(8) => dataout_from_mem(8), 
                           dataout_from_mem(7) => dataout_from_mem(7), 
                           dataout_from_mem(6) => dataout_from_mem(6), 
                           dataout_from_mem(5) => dataout_from_mem(5), 
                           dataout_from_mem(4) => dataout_from_mem(4), 
                           dataout_from_mem(3) => dataout_from_mem(3), 
                           dataout_from_mem(2) => dataout_from_mem(2), 
                           dataout_from_mem(1) => dataout_from_mem(1), 
                           dataout_from_mem(0) => dataout_from_mem(0), 
                           addr_mem(31) => addr_mem(31), addr_mem(30) => 
                           addr_mem(30), addr_mem(29) => addr_mem(29), 
                           addr_mem(28) => addr_mem(28), addr_mem(27) => 
                           addr_mem(27), addr_mem(26) => addr_mem(26), 
                           addr_mem(25) => addr_mem(25), addr_mem(24) => 
                           addr_mem(24), addr_mem(23) => addr_mem(23), 
                           addr_mem(22) => addr_mem(22), addr_mem(21) => 
                           addr_mem(21), addr_mem(20) => addr_mem(20), 
                           addr_mem(19) => addr_mem(19), addr_mem(18) => 
                           addr_mem(18), addr_mem(17) => addr_mem(17), 
                           addr_mem(16) => addr_mem(16), addr_mem(15) => 
                           addr_mem(15), addr_mem(14) => addr_mem(14), 
                           addr_mem(13) => addr_mem(13), addr_mem(12) => 
                           addr_mem(12), addr_mem(11) => addr_mem(11), 
                           addr_mem(10) => addr_mem(10), addr_mem(9) => 
                           addr_mem(9), addr_mem(8) => addr_mem(8), addr_mem(7)
                           => addr_mem(7), addr_mem(6) => addr_mem(6), 
                           addr_mem(5) => addr_mem(5), addr_mem(4) => 
                           addr_mem(4), addr_mem(3) => addr_mem(3), addr_mem(2)
                           => addr_mem(2), addr_mem(1) => addr_mem(1), 
                           addr_mem(0) => addr_mem(0), datain_mem(31) => 
                           datain_mem(31), datain_mem(30) => datain_mem(30), 
                           datain_mem(29) => datain_mem(29), datain_mem(28) => 
                           datain_mem(28), datain_mem(27) => datain_mem(27), 
                           datain_mem(26) => datain_mem(26), datain_mem(25) => 
                           datain_mem(25), datain_mem(24) => datain_mem(24), 
                           datain_mem(23) => datain_mem(23), datain_mem(22) => 
                           datain_mem(22), datain_mem(21) => datain_mem(21), 
                           datain_mem(20) => datain_mem(20), datain_mem(19) => 
                           datain_mem(19), datain_mem(18) => datain_mem(18), 
                           datain_mem(17) => datain_mem(17), datain_mem(16) => 
                           datain_mem(16), datain_mem(15) => datain_mem(15), 
                           datain_mem(14) => datain_mem(14), datain_mem(13) => 
                           datain_mem(13), datain_mem(12) => datain_mem(12), 
                           datain_mem(11) => datain_mem(11), datain_mem(10) => 
                           datain_mem(10), datain_mem(9) => datain_mem(9), 
                           datain_mem(8) => datain_mem(8), datain_mem(7) => 
                           datain_mem(7), datain_mem(6) => datain_mem(6), 
                           datain_mem(5) => datain_mem(5), datain_mem(4) => 
                           datain_mem(4), datain_mem(3) => datain_mem(3), 
                           datain_mem(2) => datain_mem(2), datain_mem(1) => 
                           datain_mem(1), datain_mem(0) => datain_mem(0), 
                           b_op_mem => b_op_mem_i, j_op_mem => j_op_mem_i, 
                           jal_op_mem => jal_op_mem_i, MemtoReg_wb => 
                           MemtoReg_wb_i, pipe_out(31) => dlx_data_out(31), 
                           pipe_out(30) => dlx_data_out(30), pipe_out(29) => 
                           dlx_data_out(29), pipe_out(28) => dlx_data_out(28), 
                           pipe_out(27) => dlx_data_out(27), pipe_out(26) => 
                           dlx_data_out(26), pipe_out(25) => dlx_data_out(25), 
                           pipe_out(24) => dlx_data_out(24), pipe_out(23) => 
                           dlx_data_out(23), pipe_out(22) => dlx_data_out(22), 
                           pipe_out(21) => dlx_data_out(21), pipe_out(20) => 
                           dlx_data_out(20), pipe_out(19) => dlx_data_out(19), 
                           pipe_out(18) => dlx_data_out(18), pipe_out(17) => 
                           dlx_data_out(17), pipe_out(16) => dlx_data_out(16), 
                           pipe_out(15) => dlx_data_out(15), pipe_out(14) => 
                           dlx_data_out(14), pipe_out(13) => dlx_data_out(13), 
                           pipe_out(12) => dlx_data_out(12), pipe_out(11) => 
                           dlx_data_out(11), pipe_out(10) => dlx_data_out(10), 
                           pipe_out(9) => dlx_data_out(9), pipe_out(8) => 
                           dlx_data_out(8), pipe_out(7) => dlx_data_out(7), 
                           pipe_out(6) => dlx_data_out(6), pipe_out(5) => 
                           dlx_data_out(5), pipe_out(4) => dlx_data_out(4), 
                           pipe_out(3) => dlx_data_out(3), pipe_out(2) => 
                           dlx_data_out(2), pipe_out(1) => dlx_data_out(1), 
                           pipe_out(0) => dlx_data_out(0));
   FF1_en : flip_flop_0 port map( D => n4, CK => Clk, Enable_n => X_Logic0_port
                           , RESET_n => X_Logic1_port, Q => CU_en1);
   FF2_en : flip_flop_1 port map( D => CU_en1, CK => Clk, Enable_n => 
                           X_Logic0_port, RESET_n => X_Logic1_port, Q => CU_en2
                           );
   CU_I : 
                           dlx_cu_MICROCODE_MEM_SIZE45_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 
                           port map( Clk => Clk, Rst => Rst, En => CU_en2, 
                           IR_opcode(5) => Opcode_i_5_port, IR_opcode(4) => 
                           Opcode_i_4_port, IR_opcode(3) => Opcode_i_3_port, 
                           IR_opcode(2) => Opcode_i_2_port, IR_opcode(1) => 
                           Opcode_i_1_port, IR_opcode(0) => Opcode_i_0_port, 
                           IR_func(10) => Func_i_10_port, IR_func(9) => 
                           Func_i_9_port, IR_func(8) => Func_i_8_port, 
                           IR_func(7) => Func_i_7_port, IR_func(6) => 
                           Func_i_6_port, IR_func(5) => Func_i_5_port, 
                           IR_func(4) => Func_i_4_port, IR_func(3) => 
                           Func_i_3_port, IR_func(2) => Func_i_2_port, 
                           IR_func(1) => Func_i_1_port, IR_func(0) => 
                           Func_i_0_port, PC_OP => n_1272, EN_REG_IF => 
                           en_reg_if_i, EN_REG_ID => en_reg_id_i, RD1 => RD1_i,
                           RD2 => RD2_i, SEL_EX => n_1273, EN_REG_EX => 
                           en_reg_ex_i, SEL_MUX_RW => n_1274, ALU_OPCODE(3) => 
                           alu_sel_i_3_port, ALU_OPCODE(2) => alu_sel_i_2_port,
                           ALU_OPCODE(1) => alu_sel_i_1_port, ALU_OPCODE(0) => 
                           alu_sel_i_0_port, EN_REG_MEM => en_reg_mem_i, 
                           MEM_EN_MEM => MEM_EN_MEM, RD_MEM => n_1275, WR_MEM 
                           => n_1276, B_OP_MEM => n_1277, J_OP_MEM => n_1278, 
                           JAL_OP_MEM => n_1279, MEM_TO_REG_WB => MemtoReg_wb_i
                           , WR => n_1280);
   U14 : INV_X1 port map( A => Rst, ZN => n4);

end SYN_dlx_rtl;
